ftdi_out_io_buffer_5b_inst : ftdi_out_io_buffer_5b PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
