library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.farm_rmap_mem_area_ffee_aeb_pkg.all;
use work.farm_avalon_mm_rmap_ffee_aeb_pkg.all;

entity farm_rmap_mem_area_ffee_aeb_write_ent is
	port(
		clk_i               : in  std_logic;
		rst_i               : in  std_logic;
		fee_rmap_i          : in  t_farm_ffee_aeb_rmap_write_in;
		avalon_mm_rmap_i    : in  t_farm_avalon_mm_rmap_ffee_aeb_write_in;
		fee_rmap_o          : out t_farm_ffee_aeb_rmap_write_out;
		avalon_mm_rmap_o    : out t_farm_avalon_mm_rmap_ffee_aeb_write_out;
		rmap_registers_wr_o : out t_rmap_memory_wr_area
	);
end entity farm_rmap_mem_area_ffee_aeb_write_ent;

architecture RTL of farm_rmap_mem_area_ffee_aeb_write_ent is

	signal s_data_acquired : std_logic;

begin

	p_farm_rmap_mem_area_ffee_aeb_write : process(clk_i, rst_i) is
		procedure p_ffee_aeb_reg_reset is
		begin

-- Write Registers Reset/Default State

-- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_0 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "NEW_STATE" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.new_state <= "0000";
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "SET_STATE" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.set_state <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "AEB_RESET" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.aeb_reset <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_1 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_DATA_RD" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_data_rd <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_WR" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_wr <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_RD" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_rd <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "DAC_WR" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.dac_wr <= '0';
-- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_2" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_2 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_0 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "WATCH-DOG_DIS" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.watchdog_dis <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "INT_SYNC" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.int_sync <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_1 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP_CDS_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp_cds_en <= '1';
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP2_CAL_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp2_cal_en <= '1';
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP1_CAL_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp1_cal_en <= '1';
-- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_2" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_2 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_SW" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_sw <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_0 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN3" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van3 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN2" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van2 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN1" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van1 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCLK" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vclk <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCCD" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vccd <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_VASP" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_vasp <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_1 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_PIX_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_pix_en <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_PIX_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_pix_en <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_ADC_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_adc_en <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_ADC_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_adc_en <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_RESET" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_reset <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_RESET" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_reset <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_ADC" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_adc <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_EN_P5V0" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_en_p5v0 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_EN_P5V0" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_en_p5v0 <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "PT1000_CAL_ON_N" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.pt1000_cal_on_n <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "EN_V_MUX_N" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.en_v_mux_n <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_PWDN_N" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_pwdn_n <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_PWDN_N" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_pwdn_n <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC_CLK_EN" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc_clk_en <= '0';
-- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_2" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_2 <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_CCDID" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_ccdid <= "00";
-- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_COLS" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_cols <= std_logic_vector(to_unsigned(32, 14));
-- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_ROWS" Field
rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_rows <= std_logic_vector(to_unsigned(32, 14));
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP_CFG_ADDR" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp_cfg_addr <= (others => '0');
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_CFG_DATA" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_cfg_data <= (others => '0');
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_CFG_DATA" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_cfg_data <= (others => '0');
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_SELECT" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_select <= '0';
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_SELECT" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_select <= '0';
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "CALIBRATION_START" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.calibration_start <= '0';
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_READ_START" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_read_start <= '0';
-- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_WRITE_START" Field
rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_write_start <= '0';
-- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_0 <= (others => '0');
-- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VOG" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vog <= x"800";
-- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_1 <= (others => '0');
-- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VRD" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vrd <= x"800";
-- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_0 <= (others => '0');
-- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "DAC_VOD" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.dac_vod <= x"800";
-- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_1 <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCCD_ON" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vccd_on <= x"00";
-- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCLK_ON" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vclk_on <= x"63";
-- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN1_ON" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van1_on <= x"C8";
-- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN2_ON" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van2_on <= x"C8";
-- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN3_ON" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van3_on <= x"C8";
-- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCCD_OFF" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vccd_off <= x"C8";
-- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCLK_OFF" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vclk_off <= x"63";
-- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN1_OFF" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van1_off <= x"00";
-- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN2_OFF" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van2_off <= x"00";
-- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN3_OFF" Field
rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van3_off <= x"00";
-- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved <= (others => '0');
-- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_0 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SPIRST" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.spirst <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "MUXMOD" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.muxmod <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "BYPAS" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.bypas <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CLKENB" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.clkenb <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CHOP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.chop <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "STAT" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.stat <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_1 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "IDLMOD" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.idlmod <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DLY" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.dly <= "100";
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SBCS" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.sbcs <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DRATE" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.drate <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainp <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINN" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainn <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DIFF" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.diff <= x"3F";
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain7 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain6 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain5 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain4 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain3 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain2 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain1 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain0 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN15" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain15 <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN14" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain14 <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN13" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain13 <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN12" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain12 <= '1';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN11" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain11 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN10" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain10 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN9" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain9 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN8" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain8 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "REF" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ref <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "GAIN" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.gain <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "TEMP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.temp <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "VCC" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.vcc <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_1 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "OFFSET" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.offset <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio7 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio6 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio5 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio4 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio3 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio2 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio1 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio0 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio7 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio6 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio5 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio4 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio3 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio2 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio1 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio0 <= '0';
-- AEB General Configuration Area Register "ADC1_CONFIG_3" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_0 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SPIRST" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.spirst <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "MUXMOD" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.muxmod <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "BYPAS" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.bypas <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CLKENB" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.clkenb <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CHOP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.chop <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "STAT" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.stat <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_1 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "IDLMOD" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.idlmod <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DLY" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.dly <= "100";
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SBCS" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.sbcs <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DRATE" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.drate <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainp <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINN" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainn <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DIFF" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.diff <= x"8F";
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain7 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain6 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain5 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain4 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain3 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain2 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain1 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain0 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN15" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain15 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN14" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain14 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN13" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain13 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN12" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain12 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN11" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain11 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN10" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain10 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN9" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain9 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN8" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain8 <= '1';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "REF" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ref <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "GAIN" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.gain <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "TEMP" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.temp <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "VCC" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.vcc <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_1 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "OFFSET" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.offset <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio7 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio6 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio5 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio4 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio3 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio2 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio1 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio0 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO7" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio7 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO6" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio6 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO5" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio5 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO4" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio4 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO3" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio3 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO2" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio2 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO1" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio1 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO0" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio0 <= '0';
-- AEB General Configuration Area Register "ADC2_CONFIG_3" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_CCD_ENABLE" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ccd_enable <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPARE" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_spare <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTLINE" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstline <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTFRM" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstfrm <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_VASPCLAMP" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_vaspclamp <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_PRECLAMP" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_preclamp <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IG" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ig <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TG" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tg <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_DG" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_dg <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHIR" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphir <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SW" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sw <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI3" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi3 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI2" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi2 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi1 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI4" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi4 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI3" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi3 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI2" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi2 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi1 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI4" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi4 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI3" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi3 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI2" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi2 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi1 <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_1 <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_1" : "ADC_CLK_DIV" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.adc_clk_div <= "0011111";
-- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_low_pos <= x"0E";
-- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_high_pos <= x"1F";
-- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_high_pos <= x"11";
-- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_high_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_high_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_high_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_high_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_LOW_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_low_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_HIGH_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_high_pos <= x"00";
-- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_CTRL" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_ctrl <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_5" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.reserved <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_EN_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_en_pos <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_CTRL_INV" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_ctrl_inv <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_0 <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_DIS_POS" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_dis_pos <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_1 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_9" : "FT_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.ft_loop_cnt <= "00100011000101";
-- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_ENABLED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_enabled <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_1 <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_loop_cnt <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_ENABLED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_enabled <= '1';
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_0 <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_loop_cnt <= "00100011000101";
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_ENABLED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_enabled <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_1 <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_loop_cnt <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_ENABLED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_enabled <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_11" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.reserved <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_loop_cnt <= "00101000000000";
-- AEB General Configuration Area Register "SEQ_CONFIG_11" : "PIX_LOOP_CNT_WORD_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.pix_loop_cnt_word_1 <= x"0000";
-- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PIX_LOOP_CNT_WORD_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pix_loop_cnt_word_0 <= x"08C5";
-- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_ENABLED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_enabled <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_12" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.reserved <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_loop_cnt <= "01000110001010";
-- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT1_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int1_loop_cnt <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_1 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT2_LOOP_CNT" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int2_loop_cnt <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_0" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_0 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_14" : "SPHI_INV" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.sphi_inv <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_1" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_1 <= (others => '0');
-- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RPHI_INV" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.rphi_inv <= '0';
-- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_2" Field
rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_2 <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved <= (others => '0');
-- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved <= (others => '0');
-- AEB Housekeeping Area Register "AEB_STATUS" : "AEB_STATUS" Field
rmap_registers_wr_o.aeb_hk_aeb_status.aeb_status <= (others => '0');
-- AEB Housekeeping Area Register "AEB_STATUS" : "VASP2_CFG_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.vasp2_cfg_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "VASP1_CFG_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.vasp1_cfg_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "DAC_CFG_WR_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.dac_cfg_wr_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_RD_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_rd_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_WR_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_wr_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_DAT_RD_RUN" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_dat_rd_run <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_ERROR" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_error <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC2_LU" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc2_lu <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC1_LU" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc1_lu <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_DAT_RD" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_dat_rd <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_RD" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_rd <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_WR" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_wr <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC2_BUSY" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc2_busy <= '0';
-- AEB Housekeeping Area Register "AEB_STATUS" : "ADC1_BUSY" Field
rmap_registers_wr_o.aeb_hk_aeb_status.adc1_busy <= '0';
-- AEB Housekeeping Area Register "TIMESTAMP_1" : "TIMESTAMP_DWORD_1" Field
rmap_registers_wr_o.aeb_hk_timestamp_1.timestamp_dword_1 <= (others => '0');
-- AEB Housekeeping Area Register "TIMESTAMP_2" : "TIMESTAMP_DWORD_0" Field
rmap_registers_wr_o.aeb_hk_timestamp_2.timestamp_dword_0 <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "ADC_CHX_DATA_T_VASP_L" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.adc_chx_data_t_vasp_l <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "ADC_CHX_DATA_T_VASP_R" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.adc_chx_data_t_vasp_r <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "ADC_CHX_DATA_T_BIAS_P" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.adc_chx_data_t_bias_p <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "ADC_CHX_DATA_T_HK_P" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.adc_chx_data_t_hk_p <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "ADC_CHX_DATA_T_TOU_1_P" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.adc_chx_data_t_tou_1_p <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "ADC_CHX_DATA_T_TOU_2_P" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.adc_chx_data_t_tou_2_p <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "ADC_CHX_DATA_HK_VODE" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.adc_chx_data_hk_vode <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "ADC_CHX_DATA_HK_VODF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.adc_chx_data_hk_vodf <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "ADC_CHX_DATA_HK_VRD" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.adc_chx_data_hk_vrd <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "ADC_CHX_DATA_HK_VOG" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.adc_chx_data_hk_vog <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "ADC_CHX_DATA_T_CCD" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.adc_chx_data_t_ccd <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "ADC_CHX_DATA_T_REF1K_MEA" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.adc_chx_data_t_ref1k_mea <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "ADC_CHX_DATA_T_REF649R_MEA" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.adc_chx_data_t_ref649r_mea <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "ADC_CHX_DATA_HK_ANA_N5V" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.adc_chx_data_hk_ana_n5v <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "ADC_CHX_DATA_S_REF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.adc_chx_data_s_ref <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "ADC_CHX_DATA_HK_CCD_P31V" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.adc_chx_data_hk_ccd_p31v <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "ADC_CHX_DATA_HK_CLK_P15V" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.adc_chx_data_hk_clk_p15v <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "ADC_CHX_DATA_HK_ANA_P5V" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.adc_chx_data_hk_ana_p5v <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "ADC_CHX_DATA_HK_ANA_P3V3" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.adc_chx_data_hk_ana_p3v3 <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "ADC_CHX_DATA_HK_DIG_P3V3" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.adc_chx_data_hk_dig_p3v3 <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "NEW" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.new_data <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "OVF" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.ovf <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "SUPPLY" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.supply <= '0';
-- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "CHID" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.chid <= (others => '0');
-- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "ADC_CHX_DATA_ADC_REF_BUF_2" Field
rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.adc_chx_data_adc_ref_buf_2 <= (others => '0');
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SPIRST" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.spirst <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "MUXMOD" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.muxmod <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "BYPAS" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.bypas <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "CLKENB" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.clkenb <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "CHOP" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.chop <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "STAT" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.stat <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "IDLMOD" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.idlmod <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SBCS1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.sbcs1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SBCS0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.sbcs0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DRATE1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.drate1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DRATE0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.drate0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF7" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff7 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF6" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff6 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF5" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff5 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF4" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff4 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN7" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain7 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN6" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain6 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN5" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain5 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN4" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain4 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN15" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain15 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN14" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain14 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN13" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain13 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN12" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain12 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN11" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain11 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN10" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain10 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN9" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain9 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN8" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain8 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "REF" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ref <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "GAIN" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.gain <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "TEMP" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.temp <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "VCC" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.vcc <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "OFFSET" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.offset <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO7" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio7 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO6" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio6 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO5" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio5 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO4" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio4 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio0 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO7" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio7 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO6" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio6 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO5" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio5 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO4" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio4 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO3" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio3 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO2" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio2 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO1" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio1 <= '0';
-- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO0" Field
rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SPIRST" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.spirst <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "MUXMOD" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.muxmod <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "BYPAS" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.bypas <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "CLKENB" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.clkenb <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "CHOP" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.chop <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "STAT" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.stat <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "IDLMOD" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.idlmod <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SBCS1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.sbcs1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SBCS0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.sbcs0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DRATE1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.drate1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DRATE0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.drate0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF7" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff7 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF6" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff6 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF5" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff5 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF4" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff4 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN7" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain7 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN6" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain6 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN5" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain5 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN4" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain4 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN15" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain15 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN14" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain14 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN13" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain13 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN12" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain12 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN11" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain11 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN10" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain10 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN9" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain9 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN8" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain8 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "REF" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ref <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "GAIN" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.gain <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "TEMP" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.temp <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "VCC" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.vcc <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "OFFSET" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.offset <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO7" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio7 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO6" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio6 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO5" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio5 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO4" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio4 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio0 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO7" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio7 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO6" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio6 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO5" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio5 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO4" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio4 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO3" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio3 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO2" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio2 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO1" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio1 <= '0';
-- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO0" Field
rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio0 <= '0';
-- AEB Housekeeping Area Register "VASP_RD_CONFIG" : "VASP1_READ_DATA" Field
rmap_registers_wr_o.aeb_hk_vasp_rd_config.vasp1_read_data <= (others => '0');
-- AEB Housekeeping Area Register "VASP_RD_CONFIG" : "VASP2_READ_DATA" Field
rmap_registers_wr_o.aeb_hk_vasp_rd_config.vasp2_read_data <= (others => '0');
-- AEB Housekeeping Area Register "REVISION_ID_1" : "FPGA_VERSION" Field
rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_version <= (others => '0');
-- AEB Housekeeping Area Register "REVISION_ID_1" : "FPGA_DATE" Field
rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_date <= (others => '0');
-- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_TIME_H" Field
rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_time_h <= (others => '0');
-- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_TIME_M" Field
rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_time_m <= (others => '0');
-- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_SVN" Field
rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_svn <= (others => '0');

		end procedure p_ffee_aeb_reg_reset;

		procedure p_ffee_aeb_reg_trigger is
		begin

-- Write Registers Triggers Reset


		end procedure p_ffee_aeb_reg_trigger;

		procedure p_ffee_aeb_mem_wr(wr_addr_i : std_logic_vector) is
		begin

-- MemArea Write Data
case (wr_addr_i(31 downto 0)) is
  -- Case for access to all memory area

  when (x"00000000") =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "AEB_RESET" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.aeb_reset <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "SET_STATE" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.set_state <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "NEW_STATE" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.new_state <= fee_rmap_i.writedata(5 downto 2);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000001") =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "DAC_WR" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.dac_wr <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_RD" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_rd <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_WR" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_wr <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_DATA_RD" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_data_rd <= fee_rmap_i.writedata(3);
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_1 <= fee_rmap_i.writedata(7 downto 4);

  when (x"00000002") =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_2(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000003") =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_2(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000004") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "INT_SYNC" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.int_sync <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "WATCH-DOG_DIS" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.watchdog_dis <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_0 <= fee_rmap_i.writedata(7 downto 2);

  when (x"00000005") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP1_CAL_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp1_cal_en <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP2_CAL_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp2_cal_en <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP_CDS_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp_cds_en <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_1 <= fee_rmap_i.writedata(7 downto 3);

  when (x"00000006") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_2(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000007") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_2(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000008") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000009") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000000A") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000000B") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000000C") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCCD" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vccd <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCLK" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vclk <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN1" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van1 <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van2 <= fee_rmap_i.writedata(3);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN3" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van3 <= fee_rmap_i.writedata(4);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_0 <= fee_rmap_i.writedata(6 downto 5);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_SW" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_sw <= fee_rmap_i.writedata(7);

  when (x"0000000D") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_RESET" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_reset <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_RESET" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_reset <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_ADC_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_adc_en <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_ADC_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_adc_en <= fee_rmap_i.writedata(3);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_PIX_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_pix_en <= fee_rmap_i.writedata(4);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_PIX_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_pix_en <= fee_rmap_i.writedata(5);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_1 <= fee_rmap_i.writedata(6);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_VASP" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_vasp <= fee_rmap_i.writedata(7);

  when (x"0000000E") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC_CLK_EN" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc_clk_en <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_PWDN_N" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_pwdn_n <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_PWDN_N" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_pwdn_n <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "EN_V_MUX_N" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.en_v_mux_n <= fee_rmap_i.writedata(3);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "PT1000_CAL_ON_N" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.pt1000_cal_on_n <= fee_rmap_i.writedata(4);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_EN_P5V0" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_en_p5v0 <= fee_rmap_i.writedata(5);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_EN_P5V0" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_en_p5v0 <= fee_rmap_i.writedata(6);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_ADC" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_adc <= fee_rmap_i.writedata(7);

  when (x"0000000F") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_2 <= fee_rmap_i.writedata;

  when (x"00000010") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_COLS" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_cols(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_CCDID" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_ccdid <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000011") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_COLS" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_cols(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000012") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_ROWS" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_rows(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.reserved <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000013") =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_ROWS" Field
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_rows(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000014") =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP_CFG_ADDR" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp_cfg_addr <= fee_rmap_i.writedata;

  when (x"00000015") =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_CFG_DATA" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_cfg_data <= fee_rmap_i.writedata;

  when (x"00000016") =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_CFG_DATA" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_cfg_data <= fee_rmap_i.writedata;

  when (x"00000017") =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_WRITE_START" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_write_start <= fee_rmap_i.writedata(0);
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_READ_START" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_read_start <= fee_rmap_i.writedata(1);
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "CALIBRATION_START" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.calibration_start <= fee_rmap_i.writedata(2);
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_SELECT" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_select <= fee_rmap_i.writedata(3);
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_SELECT" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_select <= fee_rmap_i.writedata(4);
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.reserved <= fee_rmap_i.writedata(7 downto 5);

  when (x"00000018") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VOG" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vog(11 downto 8) <= fee_rmap_i.writedata(3 downto 0);
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_0 <= fee_rmap_i.writedata(7 downto 4);

  when (x"00000019") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VOG" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vog(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000001A") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VRD" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vrd(11 downto 8) <= fee_rmap_i.writedata(3 downto 0);
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_1 <= fee_rmap_i.writedata(7 downto 4);

  when (x"0000001B") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VRD" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vrd(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000001C") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "DAC_VOD" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.dac_vod(11 downto 8) <= fee_rmap_i.writedata(3 downto 0);
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_0 <= fee_rmap_i.writedata(7 downto 4);

  when (x"0000001D") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "DAC_VOD" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.dac_vod(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000001E") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_1(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000001F") =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_1(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000020") =>
      -- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000021") =>
      -- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000022") =>
      -- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000023") =>
      -- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000024") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCCD_ON" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vccd_on <= fee_rmap_i.writedata;

  when (x"00000025") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCLK_ON" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vclk_on <= fee_rmap_i.writedata;

  when (x"00000026") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN1_ON" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van1_on <= fee_rmap_i.writedata;

  when (x"00000027") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN2_ON" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van2_on <= fee_rmap_i.writedata;

  when (x"00000028") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN3_ON" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van3_on <= fee_rmap_i.writedata;

  when (x"00000029") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCCD_OFF" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vccd_off <= fee_rmap_i.writedata;

  when (x"0000002A") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCLK_OFF" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vclk_off <= fee_rmap_i.writedata;

  when (x"0000002B") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN1_OFF" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van1_off <= fee_rmap_i.writedata;

  when (x"0000002C") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN2_OFF" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van2_off <= fee_rmap_i.writedata;

  when (x"0000002D") =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN3_OFF" Field
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van3_off <= fee_rmap_i.writedata;

  when (x"00000030") =>
      -- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000031") =>
      -- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000032") =>
      -- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000033") =>
      -- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000034") =>
      -- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000035") =>
      -- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000036") =>
      -- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000037") =>
      -- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000038") =>
      -- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000039") =>
      -- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000003A") =>
      -- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000003B") =>
      -- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000003C") =>
      -- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000003D") =>
      -- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000003E") =>
      -- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000003F") =>
      -- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000040") =>
      -- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000041") =>
      -- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000042") =>
      -- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000043") =>
      -- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000044") =>
      -- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000045") =>
      -- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000046") =>
      -- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000047") =>
      -- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000048") =>
      -- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000049") =>
      -- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000004A") =>
      -- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000004B") =>
      -- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000004C") =>
      -- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000004D") =>
      -- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000004E") =>
      -- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000004F") =>
      -- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000050") =>
      -- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000051") =>
      -- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000052") =>
      -- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000053") =>
      -- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000054") =>
      -- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000055") =>
      -- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000056") =>
      -- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000057") =>
      -- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000058") =>
      -- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000059") =>
      -- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000005A") =>
      -- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000005B") =>
      -- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000005C") =>
      -- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000005D") =>
      -- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000005E") =>
      -- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000005F") =>
      -- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000060") =>
      -- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000061") =>
      -- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000062") =>
      -- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000063") =>
      -- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000064") =>
      -- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000065") =>
      -- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000066") =>
      -- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000067") =>
      -- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000068") =>
      -- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000069") =>
      -- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000006A") =>
      -- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000006B") =>
      -- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000006C") =>
      -- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000006D") =>
      -- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000006E") =>
      -- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000006F") =>
      -- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000070") =>
      -- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000071") =>
      -- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000072") =>
      -- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000073") =>
      -- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000074") =>
      -- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000075") =>
      -- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000076") =>
      -- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000077") =>
      -- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000078") =>
      -- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000079") =>
      -- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000007A") =>
      -- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000007B") =>
      -- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000007C") =>
      -- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000007D") =>
      -- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000007E") =>
      -- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000007F") =>
      -- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000080") =>
      -- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000081") =>
      -- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000082") =>
      -- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000083") =>
      -- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000084") =>
      -- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000085") =>
      -- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000086") =>
      -- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000087") =>
      -- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000088") =>
      -- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000089") =>
      -- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000008A") =>
      -- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000008B") =>
      -- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000008C") =>
      -- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000008D") =>
      -- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000008E") =>
      -- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000008F") =>
      -- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000090") =>
      -- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000091") =>
      -- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000092") =>
      -- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000093") =>
      -- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000094") =>
      -- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000095") =>
      -- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000096") =>
      -- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000097") =>
      -- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000098") =>
      -- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000099") =>
      -- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000009A") =>
      -- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000009B") =>
      -- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000009C") =>
      -- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000009D") =>
      -- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000009E") =>
      -- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000009F") =>
      -- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000A0") =>
      -- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000A1") =>
      -- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000A2") =>
      -- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000A3") =>
      -- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000A4") =>
      -- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000A5") =>
      -- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000A6") =>
      -- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000A7") =>
      -- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000A8") =>
      -- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000A9") =>
      -- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000AA") =>
      -- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000AB") =>
      -- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000AC") =>
      -- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000AD") =>
      -- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000AE") =>
      -- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000AF") =>
      -- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000B0") =>
      -- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000B1") =>
      -- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000B2") =>
      -- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000B3") =>
      -- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000B4") =>
      -- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000B5") =>
      -- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000B6") =>
      -- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000B7") =>
      -- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000B8") =>
      -- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000B9") =>
      -- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000BA") =>
      -- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000BB") =>
      -- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000BC") =>
      -- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000BD") =>
      -- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000BE") =>
      -- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000BF") =>
      -- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000C0") =>
      -- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000C1") =>
      -- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000C2") =>
      -- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000C3") =>
      -- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000C4") =>
      -- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000C5") =>
      -- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000C6") =>
      -- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000C7") =>
      -- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000C8") =>
      -- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000C9") =>
      -- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000CA") =>
      -- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000CB") =>
      -- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000CC") =>
      -- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000CD") =>
      -- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000CE") =>
      -- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000CF") =>
      -- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000D0") =>
      -- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000D1") =>
      -- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000D2") =>
      -- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000D3") =>
      -- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000D4") =>
      -- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000D5") =>
      -- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000D6") =>
      -- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000D7") =>
      -- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000D8") =>
      -- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000D9") =>
      -- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000DA") =>
      -- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000DB") =>
      -- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000DC") =>
      -- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000DD") =>
      -- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000DE") =>
      -- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000DF") =>
      -- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000E0") =>
      -- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000E1") =>
      -- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000E2") =>
      -- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000E3") =>
      -- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000E4") =>
      -- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000E5") =>
      -- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000E6") =>
      -- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000E7") =>
      -- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000E8") =>
      -- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000E9") =>
      -- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000EA") =>
      -- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000EB") =>
      -- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000EC") =>
      -- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000ED") =>
      -- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000EE") =>
      -- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000EF") =>
      -- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000F0") =>
      -- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000F1") =>
      -- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000F2") =>
      -- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000F3") =>
      -- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000F4") =>
      -- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000F5") =>
      -- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000F6") =>
      -- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000F7") =>
      -- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000F8") =>
      -- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000F9") =>
      -- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000FA") =>
      -- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000FB") =>
      -- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000000FC") =>
      -- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000000FD") =>
      -- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000000FE") =>
      -- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000000FF") =>
      -- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000100") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_1 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "STAT" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.stat <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CHOP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.chop <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CLKENB" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.clkenb <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "BYPAS" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.bypas <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "MUXMOD" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.muxmod <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SPIRST" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.spirst <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_0 <= fee_rmap_i.writedata(7);

  when (x"00000101") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DRATE" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.drate <= fee_rmap_i.writedata(1 downto 0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SBCS" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.sbcs <= fee_rmap_i.writedata(3 downto 2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DLY" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.dly <= fee_rmap_i.writedata(6 downto 4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "IDLMOD" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.idlmod <= fee_rmap_i.writedata(7);

  when (x"00000102") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINN" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainn <= fee_rmap_i.writedata(3 downto 0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainp <= fee_rmap_i.writedata(7 downto 4);

  when (x"00000103") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DIFF" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.diff <= fee_rmap_i.writedata;

  when (x"00000104") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain7 <= fee_rmap_i.writedata(7);

  when (x"00000105") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN8" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain8 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN9" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain9 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN10" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain10 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN11" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain11 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN12" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain12 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN13" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain13 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN14" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain14 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN15" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain15 <= fee_rmap_i.writedata(7);

  when (x"00000106") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "OFFSET" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.offset <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "VCC" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.vcc <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "TEMP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.temp <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "GAIN" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.gain <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "REF" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ref <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000107") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio7 <= fee_rmap_i.writedata(7);

  when (x"00000108") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio7 <= fee_rmap_i.writedata(7);

  when (x"00000109") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000010A") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000010B") =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000010C") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_1 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "STAT" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.stat <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CHOP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.chop <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CLKENB" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.clkenb <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "BYPAS" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.bypas <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "MUXMOD" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.muxmod <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SPIRST" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.spirst <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_0 <= fee_rmap_i.writedata(7);

  when (x"0000010D") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DRATE" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.drate <= fee_rmap_i.writedata(1 downto 0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SBCS" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.sbcs <= fee_rmap_i.writedata(3 downto 2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DLY" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.dly <= fee_rmap_i.writedata(6 downto 4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "IDLMOD" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.idlmod <= fee_rmap_i.writedata(7);

  when (x"0000010E") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINN" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainn <= fee_rmap_i.writedata(3 downto 0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainp <= fee_rmap_i.writedata(7 downto 4);

  when (x"0000010F") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DIFF" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.diff <= fee_rmap_i.writedata;

  when (x"00000110") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain7 <= fee_rmap_i.writedata(7);

  when (x"00000111") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN8" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain8 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN9" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain9 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN10" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain10 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN11" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain11 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN12" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain12 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN13" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain13 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN14" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain14 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN15" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain15 <= fee_rmap_i.writedata(7);

  when (x"00000112") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "OFFSET" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.offset <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "VCC" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.vcc <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "TEMP" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.temp <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "GAIN" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.gain <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "REF" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ref <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000113") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio7 <= fee_rmap_i.writedata(7);

  when (x"00000114") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO0" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio0 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO1" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio1 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO2" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio2 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO3" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio3 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO4" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio4 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO5" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio5 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO6" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio6 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO7" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio7 <= fee_rmap_i.writedata(7);

  when (x"00000115") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000116") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000117") =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000118") =>
      -- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000119") =>
      -- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000011A") =>
      -- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000011B") =>
      -- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000011C") =>
      -- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000011D") =>
      -- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000011E") =>
      -- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000011F") =>
      -- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000120") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_PRECLAMP" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_preclamp <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_VASPCLAMP" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_vaspclamp <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTFRM" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstfrm <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTLINE" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstline <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPARE" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_spare <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_CCD_ENABLE" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ccd_enable <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000121") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi1 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI2" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi2 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI3" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi3 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SW" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sw <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHIR" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphir <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_DG" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_dg <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TG" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tg <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IG" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ig <= fee_rmap_i.writedata(7);

  when (x"00000122") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi1 <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI2" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi2 <= fee_rmap_i.writedata(1);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI3" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi3 <= fee_rmap_i.writedata(2);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI4" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi4 <= fee_rmap_i.writedata(3);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi1 <= fee_rmap_i.writedata(4);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI2" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi2 <= fee_rmap_i.writedata(5);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI3" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi3 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI4" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi4 <= fee_rmap_i.writedata(7);

  when (x"00000123") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "ADC_CLK_DIV" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.adc_clk_div <= fee_rmap_i.writedata(6 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_1 <= fee_rmap_i.writedata(7);

  when (x"00000124") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_low_pos <= fee_rmap_i.writedata;

  when (x"00000125") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_high_pos <= fee_rmap_i.writedata;

  when (x"00000126") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_low_pos <= fee_rmap_i.writedata;

  when (x"00000127") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_high_pos <= fee_rmap_i.writedata;

  when (x"00000128") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_low_pos <= fee_rmap_i.writedata;

  when (x"00000129") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_high_pos <= fee_rmap_i.writedata;

  when (x"0000012A") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_low_pos <= fee_rmap_i.writedata;

  when (x"0000012B") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_high_pos <= fee_rmap_i.writedata;

  when (x"0000012C") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_low_pos <= fee_rmap_i.writedata;

  when (x"0000012D") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_high_pos <= fee_rmap_i.writedata;

  when (x"0000012E") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_low_pos <= fee_rmap_i.writedata;

  when (x"0000012F") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_high_pos <= fee_rmap_i.writedata;

  when (x"00000130") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_LOW_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_low_pos <= fee_rmap_i.writedata;

  when (x"00000131") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_HIGH_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_high_pos <= fee_rmap_i.writedata;

  when (x"00000132") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_EN_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_en_pos(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.reserved <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_CTRL" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_ctrl <= fee_rmap_i.writedata(7);

  when (x"00000133") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_EN_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_en_pos(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000134") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_DIS_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_dis_pos(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_0 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_CTRL_INV" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_ctrl_inv <= fee_rmap_i.writedata(7);

  when (x"00000135") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_DIS_POS" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_dis_pos(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000136") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_1(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000137") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_1(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000138") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000139") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000013A") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000013B") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000013C") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000013D") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000013E") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000013F") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000140") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "FT_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.ft_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000141") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "FT_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.ft_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000142") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_1 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_ENABLED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_enabled <= fee_rmap_i.writedata(7);

  when (x"00000143") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000144") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_0 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_ENABLED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_enabled <= fee_rmap_i.writedata(7);

  when (x"00000145") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000146") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_1 <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_ENABLED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_enabled <= fee_rmap_i.writedata(7);

  when (x"00000147") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000148") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.reserved <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_ENABLED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_enabled <= fee_rmap_i.writedata(7);

  when (x"00000149") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000014A") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "PIX_LOOP_CNT_WORD_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.pix_loop_cnt_word_1(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000014B") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "PIX_LOOP_CNT_WORD_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.pix_loop_cnt_word_1(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000014C") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PIX_LOOP_CNT_WORD_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pix_loop_cnt_word_0(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000014D") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PIX_LOOP_CNT_WORD_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pix_loop_cnt_word_0(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000014E") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.reserved <= fee_rmap_i.writedata(6);
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_ENABLED" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_enabled <= fee_rmap_i.writedata(7);

  when (x"0000014F") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000150") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT1_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int1_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_0 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000151") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT1_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int1_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000152") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT2_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int2_loop_cnt(13 downto 8) <= fee_rmap_i.writedata(5 downto 0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_1 <= fee_rmap_i.writedata(7 downto 6);

  when (x"00000153") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT2_LOOP_CNT" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int2_loop_cnt(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000154") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "SPHI_INV" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.sphi_inv <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_0" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_0 <= fee_rmap_i.writedata(7 downto 1);

  when (x"00000155") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RPHI_INV" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.rphi_inv <= fee_rmap_i.writedata(0);
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_1" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_1 <= fee_rmap_i.writedata(7 downto 1);

  when (x"00000156") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_2(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000157") =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_2" Field
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_2(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000158") =>
      -- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000159") =>
      -- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000015A") =>
      -- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000015B") =>
      -- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000015C") =>
      -- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000015D") =>
      -- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000015E") =>
      -- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000015F") =>
      -- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000160") =>
      -- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000161") =>
      -- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000162") =>
      -- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000163") =>
      -- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000164") =>
      -- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000165") =>
      -- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000166") =>
      -- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000167") =>
      -- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000168") =>
      -- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000169") =>
      -- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000016A") =>
      -- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000016B") =>
      -- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000016C") =>
      -- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000016D") =>
      -- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000016E") =>
      -- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000016F") =>
      -- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000170") =>
      -- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000171") =>
      -- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000172") =>
      -- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000173") =>
      -- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000174") =>
      -- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000175") =>
      -- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000176") =>
      -- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000177") =>
      -- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000178") =>
      -- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000179") =>
      -- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000017A") =>
      -- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000017B") =>
      -- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000017C") =>
      -- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000017D") =>
      -- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000017E") =>
      -- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000017F") =>
      -- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000180") =>
      -- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000181") =>
      -- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000182") =>
      -- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000183") =>
      -- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000184") =>
      -- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000185") =>
      -- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000186") =>
      -- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000187") =>
      -- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000188") =>
      -- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000189") =>
      -- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000018A") =>
      -- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000018B") =>
      -- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000018C") =>
      -- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000018D") =>
      -- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000018E") =>
      -- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000018F") =>
      -- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000190") =>
      -- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000191") =>
      -- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000192") =>
      -- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000193") =>
      -- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000194") =>
      -- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000195") =>
      -- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000196") =>
      -- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000197") =>
      -- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000198") =>
      -- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000199") =>
      -- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000019A") =>
      -- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000019B") =>
      -- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000019C") =>
      -- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000019D") =>
      -- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000019E") =>
      -- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000019F") =>
      -- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001A0") =>
      -- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001A1") =>
      -- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001A2") =>
      -- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001A3") =>
      -- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001A4") =>
      -- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001A5") =>
      -- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001A6") =>
      -- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001A7") =>
      -- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001A8") =>
      -- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001A9") =>
      -- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001AA") =>
      -- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001AB") =>
      -- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001AC") =>
      -- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001AD") =>
      -- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001AE") =>
      -- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001AF") =>
      -- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001B0") =>
      -- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001B1") =>
      -- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001B2") =>
      -- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001B3") =>
      -- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001B4") =>
      -- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001B5") =>
      -- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001B6") =>
      -- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001B7") =>
      -- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001B8") =>
      -- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001B9") =>
      -- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001BA") =>
      -- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001BB") =>
      -- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001BC") =>
      -- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001BD") =>
      -- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001BE") =>
      -- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001BF") =>
      -- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001C0") =>
      -- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001C1") =>
      -- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001C2") =>
      -- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001C3") =>
      -- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001C4") =>
      -- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001C5") =>
      -- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001C6") =>
      -- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001C7") =>
      -- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001C8") =>
      -- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001C9") =>
      -- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001CA") =>
      -- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001CB") =>
      -- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001CC") =>
      -- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001CD") =>
      -- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001CE") =>
      -- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001CF") =>
      -- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001D0") =>
      -- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001D1") =>
      -- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001D2") =>
      -- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001D3") =>
      -- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001D4") =>
      -- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001D5") =>
      -- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001D6") =>
      -- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001D7") =>
      -- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001D8") =>
      -- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001D9") =>
      -- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001DA") =>
      -- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001DB") =>
      -- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001DC") =>
      -- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001DD") =>
      -- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001DE") =>
      -- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001DF") =>
      -- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001E0") =>
      -- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001E1") =>
      -- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001E2") =>
      -- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001E3") =>
      -- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001E4") =>
      -- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001E5") =>
      -- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001E6") =>
      -- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001E7") =>
      -- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001E8") =>
      -- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001E9") =>
      -- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001EA") =>
      -- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001EB") =>
      -- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001EC") =>
      -- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001ED") =>
      -- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001EE") =>
      -- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001EF") =>
      -- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001F0") =>
      -- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001F1") =>
      -- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001F2") =>
      -- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001F3") =>
      -- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001F4") =>
      -- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001F5") =>
      -- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001F6") =>
      -- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001F7") =>
      -- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001F8") =>
      -- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001F9") =>
      -- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001FA") =>
      -- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001FB") =>
      -- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000001FC") =>
      -- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000001FD") =>
      -- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000001FE") =>
      -- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000001FF") =>
      -- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000200") =>
      -- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000201") =>
      -- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000202") =>
      -- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000203") =>
      -- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000204") =>
      -- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000205") =>
      -- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000206") =>
      -- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000207") =>
      -- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000208") =>
      -- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000209") =>
      -- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000020A") =>
      -- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000020B") =>
      -- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000020C") =>
      -- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000020D") =>
      -- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000020E") =>
      -- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000020F") =>
      -- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000210") =>
      -- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000211") =>
      -- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000212") =>
      -- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000213") =>
      -- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000214") =>
      -- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000215") =>
      -- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000216") =>
      -- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000217") =>
      -- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000218") =>
      -- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000219") =>
      -- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000021A") =>
      -- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000021B") =>
      -- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000021C") =>
      -- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000021D") =>
      -- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000021E") =>
      -- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000021F") =>
      -- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000220") =>
      -- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000221") =>
      -- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000222") =>
      -- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000223") =>
      -- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000224") =>
      -- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000225") =>
      -- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000226") =>
      -- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000227") =>
      -- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000228") =>
      -- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000229") =>
      -- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000022A") =>
      -- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000022B") =>
      -- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000022C") =>
      -- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000022D") =>
      -- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000022E") =>
      -- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000022F") =>
      -- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000230") =>
      -- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000231") =>
      -- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000232") =>
      -- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000233") =>
      -- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000234") =>
      -- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000235") =>
      -- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000236") =>
      -- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000237") =>
      -- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000238") =>
      -- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000239") =>
      -- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000023A") =>
      -- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000023B") =>
      -- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000023C") =>
      -- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000023D") =>
      -- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000023E") =>
      -- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000023F") =>
      -- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000240") =>
      -- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000241") =>
      -- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000242") =>
      -- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000243") =>
      -- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000244") =>
      -- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000245") =>
      -- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000246") =>
      -- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000247") =>
      -- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000248") =>
      -- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000249") =>
      -- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000024A") =>
      -- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000024B") =>
      -- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000024C") =>
      -- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000024D") =>
      -- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000024E") =>
      -- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000024F") =>
      -- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000250") =>
      -- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000251") =>
      -- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000252") =>
      -- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000253") =>
      -- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000254") =>
      -- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000255") =>
      -- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000256") =>
      -- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000257") =>
      -- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000258") =>
      -- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000259") =>
      -- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000025A") =>
      -- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000025B") =>
      -- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000025C") =>
      -- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000025D") =>
      -- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000025E") =>
      -- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000025F") =>
      -- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000260") =>
      -- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000261") =>
      -- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000262") =>
      -- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000263") =>
      -- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000264") =>
      -- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000265") =>
      -- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000266") =>
      -- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000267") =>
      -- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000268") =>
      -- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000269") =>
      -- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000026A") =>
      -- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000026B") =>
      -- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000026C") =>
      -- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000026D") =>
      -- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000026E") =>
      -- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000026F") =>
      -- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000270") =>
      -- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000271") =>
      -- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000272") =>
      -- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000273") =>
      -- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000274") =>
      -- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000275") =>
      -- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000276") =>
      -- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000277") =>
      -- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000278") =>
      -- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000279") =>
      -- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000027A") =>
      -- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000027B") =>
      -- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000027C") =>
      -- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000027D") =>
      -- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000027E") =>
      -- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000027F") =>
      -- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000280") =>
      -- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000281") =>
      -- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000282") =>
      -- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000283") =>
      -- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000284") =>
      -- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000285") =>
      -- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000286") =>
      -- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000287") =>
      -- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000288") =>
      -- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000289") =>
      -- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000028A") =>
      -- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000028B") =>
      -- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000028C") =>
      -- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000028D") =>
      -- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000028E") =>
      -- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000028F") =>
      -- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000290") =>
      -- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000291") =>
      -- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000292") =>
      -- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000293") =>
      -- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000294") =>
      -- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000295") =>
      -- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000296") =>
      -- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000297") =>
      -- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000298") =>
      -- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000299") =>
      -- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000029A") =>
      -- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000029B") =>
      -- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000029C") =>
      -- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000029D") =>
      -- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000029E") =>
      -- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000029F") =>
      -- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002A0") =>
      -- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002A1") =>
      -- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002A2") =>
      -- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002A3") =>
      -- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002A4") =>
      -- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002A5") =>
      -- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002A6") =>
      -- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002A7") =>
      -- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002A8") =>
      -- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002A9") =>
      -- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002AA") =>
      -- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002AB") =>
      -- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002AC") =>
      -- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002AD") =>
      -- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002AE") =>
      -- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002AF") =>
      -- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002B0") =>
      -- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002B1") =>
      -- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002B2") =>
      -- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002B3") =>
      -- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002B4") =>
      -- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002B5") =>
      -- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002B6") =>
      -- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002B7") =>
      -- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002B8") =>
      -- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002B9") =>
      -- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002BA") =>
      -- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002BB") =>
      -- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002BC") =>
      -- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002BD") =>
      -- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002BE") =>
      -- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002BF") =>
      -- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002C0") =>
      -- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002C1") =>
      -- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002C2") =>
      -- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002C3") =>
      -- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002C4") =>
      -- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002C5") =>
      -- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002C6") =>
      -- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002C7") =>
      -- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002C8") =>
      -- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002C9") =>
      -- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002CA") =>
      -- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002CB") =>
      -- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002CC") =>
      -- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002CD") =>
      -- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002CE") =>
      -- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002CF") =>
      -- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002D0") =>
      -- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002D1") =>
      -- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002D2") =>
      -- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002D3") =>
      -- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002D4") =>
      -- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002D5") =>
      -- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002D6") =>
      -- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002D7") =>
      -- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002D8") =>
      -- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002D9") =>
      -- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002DA") =>
      -- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002DB") =>
      -- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002DC") =>
      -- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002DD") =>
      -- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002DE") =>
      -- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002DF") =>
      -- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002E0") =>
      -- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002E1") =>
      -- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002E2") =>
      -- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002E3") =>
      -- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002E4") =>
      -- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002E5") =>
      -- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002E6") =>
      -- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002E7") =>
      -- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002E8") =>
      -- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002E9") =>
      -- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002EA") =>
      -- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002EB") =>
      -- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002EC") =>
      -- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002ED") =>
      -- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002EE") =>
      -- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002EF") =>
      -- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002F0") =>
      -- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002F1") =>
      -- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002F2") =>
      -- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002F3") =>
      -- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002F4") =>
      -- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002F5") =>
      -- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002F6") =>
      -- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002F7") =>
      -- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002F8") =>
      -- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002F9") =>
      -- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002FA") =>
      -- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002FB") =>
      -- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000002FC") =>
      -- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000002FD") =>
      -- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000002FE") =>
      -- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000002FF") =>
      -- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000300") =>
      -- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000301") =>
      -- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000302") =>
      -- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000303") =>
      -- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000304") =>
      -- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000305") =>
      -- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000306") =>
      -- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000307") =>
      -- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000308") =>
      -- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000309") =>
      -- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000030A") =>
      -- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000030B") =>
      -- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000030C") =>
      -- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000030D") =>
      -- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000030E") =>
      -- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000030F") =>
      -- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000310") =>
      -- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000311") =>
      -- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000312") =>
      -- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000313") =>
      -- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000314") =>
      -- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000315") =>
      -- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000316") =>
      -- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000317") =>
      -- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000318") =>
      -- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000319") =>
      -- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000031A") =>
      -- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000031B") =>
      -- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000031C") =>
      -- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000031D") =>
      -- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000031E") =>
      -- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000031F") =>
      -- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000320") =>
      -- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000321") =>
      -- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000322") =>
      -- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000323") =>
      -- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000324") =>
      -- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000325") =>
      -- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000326") =>
      -- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000327") =>
      -- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000328") =>
      -- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000329") =>
      -- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000032A") =>
      -- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000032B") =>
      -- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000032C") =>
      -- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000032D") =>
      -- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000032E") =>
      -- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000032F") =>
      -- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000330") =>
      -- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000331") =>
      -- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000332") =>
      -- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000333") =>
      -- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000334") =>
      -- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000335") =>
      -- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000336") =>
      -- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000337") =>
      -- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000338") =>
      -- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000339") =>
      -- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000033A") =>
      -- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000033B") =>
      -- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000033C") =>
      -- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000033D") =>
      -- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000033E") =>
      -- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000033F") =>
      -- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000340") =>
      -- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000341") =>
      -- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000342") =>
      -- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000343") =>
      -- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000344") =>
      -- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000345") =>
      -- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000346") =>
      -- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000347") =>
      -- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000348") =>
      -- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000349") =>
      -- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000034A") =>
      -- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000034B") =>
      -- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000034C") =>
      -- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000034D") =>
      -- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000034E") =>
      -- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000034F") =>
      -- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000350") =>
      -- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000351") =>
      -- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000352") =>
      -- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000353") =>
      -- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000354") =>
      -- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000355") =>
      -- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000356") =>
      -- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000357") =>
      -- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000358") =>
      -- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000359") =>
      -- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000035A") =>
      -- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000035B") =>
      -- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000035C") =>
      -- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000035D") =>
      -- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000035E") =>
      -- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000035F") =>
      -- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000360") =>
      -- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000361") =>
      -- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000362") =>
      -- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000363") =>
      -- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000364") =>
      -- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000365") =>
      -- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000366") =>
      -- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000367") =>
      -- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000368") =>
      -- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000369") =>
      -- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000036A") =>
      -- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000036B") =>
      -- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000036C") =>
      -- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000036D") =>
      -- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000036E") =>
      -- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000036F") =>
      -- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000370") =>
      -- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000371") =>
      -- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000372") =>
      -- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000373") =>
      -- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000374") =>
      -- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000375") =>
      -- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000376") =>
      -- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000377") =>
      -- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000378") =>
      -- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000379") =>
      -- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000037A") =>
      -- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000037B") =>
      -- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000037C") =>
      -- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000037D") =>
      -- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000037E") =>
      -- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000037F") =>
      -- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000380") =>
      -- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000381") =>
      -- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000382") =>
      -- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000383") =>
      -- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000384") =>
      -- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000385") =>
      -- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000386") =>
      -- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000387") =>
      -- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000388") =>
      -- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000389") =>
      -- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000038A") =>
      -- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000038B") =>
      -- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000038C") =>
      -- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000038D") =>
      -- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000038E") =>
      -- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000038F") =>
      -- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000390") =>
      -- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000391") =>
      -- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000392") =>
      -- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000393") =>
      -- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000394") =>
      -- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000395") =>
      -- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000396") =>
      -- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000397") =>
      -- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000398") =>
      -- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000399") =>
      -- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000039A") =>
      -- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000039B") =>
      -- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000039C") =>
      -- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000039D") =>
      -- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000039E") =>
      -- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000039F") =>
      -- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003A0") =>
      -- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003A1") =>
      -- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003A2") =>
      -- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003A3") =>
      -- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003A4") =>
      -- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003A5") =>
      -- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003A6") =>
      -- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003A7") =>
      -- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003A8") =>
      -- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003A9") =>
      -- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003AA") =>
      -- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003AB") =>
      -- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003AC") =>
      -- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003AD") =>
      -- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003AE") =>
      -- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003AF") =>
      -- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003B0") =>
      -- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003B1") =>
      -- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003B2") =>
      -- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003B3") =>
      -- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003B4") =>
      -- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003B5") =>
      -- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003B6") =>
      -- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003B7") =>
      -- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003B8") =>
      -- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003B9") =>
      -- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003BA") =>
      -- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003BB") =>
      -- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003BC") =>
      -- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003BD") =>
      -- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003BE") =>
      -- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003BF") =>
      -- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003C0") =>
      -- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003C1") =>
      -- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003C2") =>
      -- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003C3") =>
      -- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003C4") =>
      -- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003C5") =>
      -- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003C6") =>
      -- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003C7") =>
      -- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003C8") =>
      -- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003C9") =>
      -- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003CA") =>
      -- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003CB") =>
      -- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003CC") =>
      -- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003CD") =>
      -- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003CE") =>
      -- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003CF") =>
      -- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003D0") =>
      -- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003D1") =>
      -- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003D2") =>
      -- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003D3") =>
      -- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003D4") =>
      -- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003D5") =>
      -- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003D6") =>
      -- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003D7") =>
      -- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003D8") =>
      -- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003D9") =>
      -- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003DA") =>
      -- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003DB") =>
      -- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003DC") =>
      -- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003DD") =>
      -- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003DE") =>
      -- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003DF") =>
      -- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003E0") =>
      -- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003E1") =>
      -- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003E2") =>
      -- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003E3") =>
      -- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003E4") =>
      -- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003E5") =>
      -- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003E6") =>
      -- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003E7") =>
      -- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003E8") =>
      -- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003E9") =>
      -- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003EA") =>
      -- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003EB") =>
      -- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003EC") =>
      -- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003ED") =>
      -- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003EE") =>
      -- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003EF") =>
      -- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003F0") =>
      -- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003F1") =>
      -- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003F2") =>
      -- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003F3") =>
      -- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003F4") =>
      -- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003F5") =>
      -- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003F6") =>
      -- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003F7") =>
      -- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003F8") =>
      -- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003F9") =>
      -- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003FA") =>
      -- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003FB") =>
      -- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000003FC") =>
      -- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000003FD") =>
      -- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000003FE") =>
      -- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000003FF") =>
      -- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000400") =>
      -- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000401") =>
      -- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000402") =>
      -- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000403") =>
      -- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000404") =>
      -- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000405") =>
      -- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000406") =>
      -- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000407") =>
      -- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000408") =>
      -- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000409") =>
      -- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000040A") =>
      -- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000040B") =>
      -- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000040C") =>
      -- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000040D") =>
      -- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000040E") =>
      -- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000040F") =>
      -- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000410") =>
      -- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000411") =>
      -- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000412") =>
      -- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000413") =>
      -- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000414") =>
      -- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000415") =>
      -- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000416") =>
      -- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000417") =>
      -- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000418") =>
      -- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000419") =>
      -- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000041A") =>
      -- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000041B") =>
      -- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000041C") =>
      -- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000041D") =>
      -- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000041E") =>
      -- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000041F") =>
      -- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000420") =>
      -- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000421") =>
      -- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000422") =>
      -- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000423") =>
      -- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000424") =>
      -- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000425") =>
      -- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000426") =>
      -- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000427") =>
      -- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000428") =>
      -- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000429") =>
      -- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000042A") =>
      -- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000042B") =>
      -- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000042C") =>
      -- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000042D") =>
      -- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000042E") =>
      -- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000042F") =>
      -- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000430") =>
      -- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000431") =>
      -- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000432") =>
      -- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000433") =>
      -- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000434") =>
      -- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000435") =>
      -- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000436") =>
      -- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000437") =>
      -- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000438") =>
      -- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000439") =>
      -- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000043A") =>
      -- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000043B") =>
      -- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000043C") =>
      -- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000043D") =>
      -- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000043E") =>
      -- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000043F") =>
      -- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000440") =>
      -- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000441") =>
      -- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000442") =>
      -- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000443") =>
      -- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000444") =>
      -- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000445") =>
      -- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000446") =>
      -- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000447") =>
      -- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000448") =>
      -- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000449") =>
      -- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000044A") =>
      -- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000044B") =>
      -- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000044C") =>
      -- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000044D") =>
      -- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000044E") =>
      -- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000044F") =>
      -- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000450") =>
      -- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000451") =>
      -- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000452") =>
      -- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000453") =>
      -- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000454") =>
      -- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000455") =>
      -- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000456") =>
      -- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000457") =>
      -- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000458") =>
      -- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000459") =>
      -- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000045A") =>
      -- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000045B") =>
      -- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000045C") =>
      -- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000045D") =>
      -- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000045E") =>
      -- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000045F") =>
      -- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000460") =>
      -- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000461") =>
      -- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000462") =>
      -- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000463") =>
      -- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000464") =>
      -- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000465") =>
      -- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000466") =>
      -- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000467") =>
      -- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000468") =>
      -- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000469") =>
      -- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000046A") =>
      -- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000046B") =>
      -- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000046C") =>
      -- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000046D") =>
      -- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000046E") =>
      -- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000046F") =>
      -- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000470") =>
      -- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000471") =>
      -- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000472") =>
      -- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000473") =>
      -- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000474") =>
      -- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000475") =>
      -- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000476") =>
      -- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000477") =>
      -- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000478") =>
      -- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000479") =>
      -- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000047A") =>
      -- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000047B") =>
      -- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000047C") =>
      -- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000047D") =>
      -- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000047E") =>
      -- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000047F") =>
      -- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000480") =>
      -- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000481") =>
      -- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000482") =>
      -- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000483") =>
      -- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000484") =>
      -- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000485") =>
      -- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000486") =>
      -- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000487") =>
      -- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000488") =>
      -- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000489") =>
      -- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000048A") =>
      -- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000048B") =>
      -- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000048C") =>
      -- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000048D") =>
      -- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000048E") =>
      -- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000048F") =>
      -- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000490") =>
      -- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000491") =>
      -- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000492") =>
      -- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000493") =>
      -- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000494") =>
      -- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000495") =>
      -- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000496") =>
      -- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000497") =>
      -- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000498") =>
      -- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000499") =>
      -- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000049A") =>
      -- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000049B") =>
      -- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000049C") =>
      -- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000049D") =>
      -- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000049E") =>
      -- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000049F") =>
      -- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004A0") =>
      -- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004A1") =>
      -- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004A2") =>
      -- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004A3") =>
      -- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004A4") =>
      -- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004A5") =>
      -- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004A6") =>
      -- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004A7") =>
      -- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004A8") =>
      -- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004A9") =>
      -- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004AA") =>
      -- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004AB") =>
      -- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004AC") =>
      -- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004AD") =>
      -- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004AE") =>
      -- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004AF") =>
      -- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004B0") =>
      -- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004B1") =>
      -- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004B2") =>
      -- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004B3") =>
      -- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004B4") =>
      -- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004B5") =>
      -- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004B6") =>
      -- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004B7") =>
      -- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004B8") =>
      -- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004B9") =>
      -- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004BA") =>
      -- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004BB") =>
      -- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004BC") =>
      -- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004BD") =>
      -- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004BE") =>
      -- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004BF") =>
      -- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004C0") =>
      -- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004C1") =>
      -- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004C2") =>
      -- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004C3") =>
      -- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004C4") =>
      -- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004C5") =>
      -- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004C6") =>
      -- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004C7") =>
      -- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004C8") =>
      -- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004C9") =>
      -- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004CA") =>
      -- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004CB") =>
      -- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004CC") =>
      -- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004CD") =>
      -- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004CE") =>
      -- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004CF") =>
      -- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004D0") =>
      -- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004D1") =>
      -- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004D2") =>
      -- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004D3") =>
      -- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004D4") =>
      -- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004D5") =>
      -- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004D6") =>
      -- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004D7") =>
      -- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004D8") =>
      -- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004D9") =>
      -- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004DA") =>
      -- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004DB") =>
      -- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004DC") =>
      -- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004DD") =>
      -- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004DE") =>
      -- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004DF") =>
      -- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004E0") =>
      -- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004E1") =>
      -- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004E2") =>
      -- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004E3") =>
      -- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004E4") =>
      -- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004E5") =>
      -- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004E6") =>
      -- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004E7") =>
      -- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004E8") =>
      -- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004E9") =>
      -- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004EA") =>
      -- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004EB") =>
      -- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004EC") =>
      -- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004ED") =>
      -- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004EE") =>
      -- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004EF") =>
      -- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004F0") =>
      -- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004F1") =>
      -- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004F2") =>
      -- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004F3") =>
      -- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004F4") =>
      -- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004F5") =>
      -- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004F6") =>
      -- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004F7") =>
      -- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004F8") =>
      -- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004F9") =>
      -- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004FA") =>
      -- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004FB") =>
      -- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000004FC") =>
      -- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000004FD") =>
      -- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000004FE") =>
      -- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000004FF") =>
      -- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000500") =>
      -- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000501") =>
      -- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000502") =>
      -- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000503") =>
      -- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000504") =>
      -- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000505") =>
      -- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000506") =>
      -- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000507") =>
      -- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000508") =>
      -- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000509") =>
      -- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000050A") =>
      -- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000050B") =>
      -- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000050C") =>
      -- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000050D") =>
      -- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000050E") =>
      -- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000050F") =>
      -- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000510") =>
      -- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000511") =>
      -- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000512") =>
      -- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000513") =>
      -- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000514") =>
      -- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000515") =>
      -- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000516") =>
      -- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000517") =>
      -- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000518") =>
      -- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000519") =>
      -- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000051A") =>
      -- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000051B") =>
      -- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000051C") =>
      -- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000051D") =>
      -- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000051E") =>
      -- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000051F") =>
      -- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000520") =>
      -- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000521") =>
      -- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000522") =>
      -- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000523") =>
      -- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000524") =>
      -- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000525") =>
      -- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000526") =>
      -- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000527") =>
      -- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000528") =>
      -- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000529") =>
      -- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000052A") =>
      -- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000052B") =>
      -- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000052C") =>
      -- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000052D") =>
      -- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000052E") =>
      -- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000052F") =>
      -- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000530") =>
      -- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000531") =>
      -- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000532") =>
      -- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000533") =>
      -- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000534") =>
      -- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000535") =>
      -- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000536") =>
      -- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000537") =>
      -- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000538") =>
      -- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000539") =>
      -- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000053A") =>
      -- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000053B") =>
      -- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000053C") =>
      -- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000053D") =>
      -- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000053E") =>
      -- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000053F") =>
      -- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000540") =>
      -- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000541") =>
      -- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000542") =>
      -- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000543") =>
      -- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000544") =>
      -- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000545") =>
      -- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000546") =>
      -- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000547") =>
      -- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000548") =>
      -- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000549") =>
      -- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000054A") =>
      -- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000054B") =>
      -- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000054C") =>
      -- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000054D") =>
      -- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000054E") =>
      -- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000054F") =>
      -- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000550") =>
      -- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000551") =>
      -- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000552") =>
      -- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000553") =>
      -- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000554") =>
      -- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000555") =>
      -- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000556") =>
      -- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000557") =>
      -- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000558") =>
      -- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000559") =>
      -- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000055A") =>
      -- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000055B") =>
      -- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000055C") =>
      -- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000055D") =>
      -- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000055E") =>
      -- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000055F") =>
      -- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000560") =>
      -- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000561") =>
      -- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000562") =>
      -- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000563") =>
      -- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000564") =>
      -- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000565") =>
      -- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000566") =>
      -- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000567") =>
      -- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000568") =>
      -- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000569") =>
      -- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000056A") =>
      -- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000056B") =>
      -- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000056C") =>
      -- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000056D") =>
      -- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000056E") =>
      -- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000056F") =>
      -- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000570") =>
      -- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000571") =>
      -- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000572") =>
      -- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000573") =>
      -- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000574") =>
      -- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000575") =>
      -- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000576") =>
      -- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000577") =>
      -- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000578") =>
      -- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000579") =>
      -- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000057A") =>
      -- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000057B") =>
      -- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000057C") =>
      -- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000057D") =>
      -- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000057E") =>
      -- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000057F") =>
      -- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000580") =>
      -- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000581") =>
      -- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000582") =>
      -- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000583") =>
      -- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000584") =>
      -- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000585") =>
      -- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000586") =>
      -- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000587") =>
      -- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000588") =>
      -- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000589") =>
      -- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000058A") =>
      -- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000058B") =>
      -- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000058C") =>
      -- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000058D") =>
      -- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000058E") =>
      -- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000058F") =>
      -- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000590") =>
      -- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000591") =>
      -- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000592") =>
      -- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000593") =>
      -- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000594") =>
      -- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000595") =>
      -- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000596") =>
      -- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000597") =>
      -- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000598") =>
      -- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000599") =>
      -- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000059A") =>
      -- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000059B") =>
      -- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000059C") =>
      -- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000059D") =>
      -- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000059E") =>
      -- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000059F") =>
      -- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005A0") =>
      -- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005A1") =>
      -- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005A2") =>
      -- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005A3") =>
      -- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005A4") =>
      -- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005A5") =>
      -- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005A6") =>
      -- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005A7") =>
      -- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005A8") =>
      -- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005A9") =>
      -- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005AA") =>
      -- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005AB") =>
      -- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005AC") =>
      -- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005AD") =>
      -- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005AE") =>
      -- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005AF") =>
      -- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005B0") =>
      -- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005B1") =>
      -- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005B2") =>
      -- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005B3") =>
      -- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005B4") =>
      -- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005B5") =>
      -- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005B6") =>
      -- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005B7") =>
      -- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005B8") =>
      -- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005B9") =>
      -- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005BA") =>
      -- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005BB") =>
      -- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005BC") =>
      -- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005BD") =>
      -- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005BE") =>
      -- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005BF") =>
      -- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005C0") =>
      -- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005C1") =>
      -- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005C2") =>
      -- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005C3") =>
      -- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005C4") =>
      -- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005C5") =>
      -- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005C6") =>
      -- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005C7") =>
      -- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005C8") =>
      -- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005C9") =>
      -- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005CA") =>
      -- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005CB") =>
      -- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005CC") =>
      -- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005CD") =>
      -- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005CE") =>
      -- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005CF") =>
      -- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005D0") =>
      -- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005D1") =>
      -- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005D2") =>
      -- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005D3") =>
      -- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005D4") =>
      -- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005D5") =>
      -- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005D6") =>
      -- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005D7") =>
      -- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005D8") =>
      -- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005D9") =>
      -- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005DA") =>
      -- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005DB") =>
      -- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005DC") =>
      -- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005DD") =>
      -- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005DE") =>
      -- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005DF") =>
      -- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005E0") =>
      -- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005E1") =>
      -- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005E2") =>
      -- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005E3") =>
      -- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005E4") =>
      -- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005E5") =>
      -- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005E6") =>
      -- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005E7") =>
      -- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005E8") =>
      -- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005E9") =>
      -- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005EA") =>
      -- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005EB") =>
      -- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005EC") =>
      -- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005ED") =>
      -- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005EE") =>
      -- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005EF") =>
      -- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005F0") =>
      -- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005F1") =>
      -- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005F2") =>
      -- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005F3") =>
      -- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005F4") =>
      -- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005F5") =>
      -- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005F6") =>
      -- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005F7") =>
      -- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005F8") =>
      -- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005F9") =>
      -- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005FA") =>
      -- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005FB") =>
      -- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000005FC") =>
      -- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000005FD") =>
      -- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000005FE") =>
      -- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000005FF") =>
      -- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000600") =>
      -- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000601") =>
      -- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000602") =>
      -- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000603") =>
      -- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000604") =>
      -- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000605") =>
      -- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000606") =>
      -- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000607") =>
      -- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000608") =>
      -- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000609") =>
      -- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000060A") =>
      -- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000060B") =>
      -- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000060C") =>
      -- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000060D") =>
      -- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000060E") =>
      -- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000060F") =>
      -- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000610") =>
      -- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000611") =>
      -- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000612") =>
      -- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000613") =>
      -- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000614") =>
      -- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000615") =>
      -- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000616") =>
      -- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000617") =>
      -- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000618") =>
      -- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000619") =>
      -- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000061A") =>
      -- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000061B") =>
      -- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000061C") =>
      -- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000061D") =>
      -- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000061E") =>
      -- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000061F") =>
      -- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000620") =>
      -- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000621") =>
      -- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000622") =>
      -- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000623") =>
      -- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000624") =>
      -- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000625") =>
      -- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000626") =>
      -- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000627") =>
      -- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000628") =>
      -- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000629") =>
      -- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000062A") =>
      -- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000062B") =>
      -- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000062C") =>
      -- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000062D") =>
      -- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000062E") =>
      -- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000062F") =>
      -- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000630") =>
      -- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000631") =>
      -- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000632") =>
      -- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000633") =>
      -- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000634") =>
      -- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000635") =>
      -- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000636") =>
      -- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000637") =>
      -- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000638") =>
      -- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000639") =>
      -- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000063A") =>
      -- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000063B") =>
      -- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000063C") =>
      -- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000063D") =>
      -- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000063E") =>
      -- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000063F") =>
      -- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000640") =>
      -- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000641") =>
      -- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000642") =>
      -- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000643") =>
      -- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000644") =>
      -- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000645") =>
      -- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000646") =>
      -- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000647") =>
      -- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000648") =>
      -- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000649") =>
      -- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000064A") =>
      -- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000064B") =>
      -- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000064C") =>
      -- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000064D") =>
      -- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000064E") =>
      -- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000064F") =>
      -- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000650") =>
      -- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000651") =>
      -- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000652") =>
      -- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000653") =>
      -- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000654") =>
      -- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000655") =>
      -- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000656") =>
      -- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000657") =>
      -- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000658") =>
      -- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000659") =>
      -- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000065A") =>
      -- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000065B") =>
      -- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000065C") =>
      -- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000065D") =>
      -- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000065E") =>
      -- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000065F") =>
      -- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000660") =>
      -- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000661") =>
      -- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000662") =>
      -- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000663") =>
      -- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000664") =>
      -- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000665") =>
      -- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000666") =>
      -- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000667") =>
      -- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000668") =>
      -- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000669") =>
      -- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000066A") =>
      -- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000066B") =>
      -- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000066C") =>
      -- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000066D") =>
      -- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000066E") =>
      -- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000066F") =>
      -- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000670") =>
      -- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000671") =>
      -- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000672") =>
      -- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000673") =>
      -- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000674") =>
      -- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000675") =>
      -- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000676") =>
      -- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000677") =>
      -- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000678") =>
      -- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000679") =>
      -- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000067A") =>
      -- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000067B") =>
      -- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000067C") =>
      -- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000067D") =>
      -- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000067E") =>
      -- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000067F") =>
      -- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000680") =>
      -- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000681") =>
      -- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000682") =>
      -- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000683") =>
      -- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000684") =>
      -- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000685") =>
      -- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000686") =>
      -- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000687") =>
      -- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000688") =>
      -- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000689") =>
      -- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000068A") =>
      -- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000068B") =>
      -- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000068C") =>
      -- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000068D") =>
      -- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000068E") =>
      -- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000068F") =>
      -- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000690") =>
      -- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000691") =>
      -- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000692") =>
      -- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000693") =>
      -- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000694") =>
      -- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000695") =>
      -- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000696") =>
      -- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000697") =>
      -- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000698") =>
      -- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000699") =>
      -- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000069A") =>
      -- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000069B") =>
      -- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000069C") =>
      -- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000069D") =>
      -- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000069E") =>
      -- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000069F") =>
      -- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006A0") =>
      -- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006A1") =>
      -- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006A2") =>
      -- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006A3") =>
      -- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006A4") =>
      -- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006A5") =>
      -- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006A6") =>
      -- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006A7") =>
      -- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006A8") =>
      -- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006A9") =>
      -- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006AA") =>
      -- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006AB") =>
      -- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006AC") =>
      -- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006AD") =>
      -- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006AE") =>
      -- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006AF") =>
      -- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006B0") =>
      -- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006B1") =>
      -- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006B2") =>
      -- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006B3") =>
      -- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006B4") =>
      -- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006B5") =>
      -- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006B6") =>
      -- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006B7") =>
      -- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006B8") =>
      -- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006B9") =>
      -- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006BA") =>
      -- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006BB") =>
      -- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006BC") =>
      -- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006BD") =>
      -- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006BE") =>
      -- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006BF") =>
      -- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006C0") =>
      -- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006C1") =>
      -- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006C2") =>
      -- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006C3") =>
      -- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006C4") =>
      -- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006C5") =>
      -- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006C6") =>
      -- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006C7") =>
      -- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006C8") =>
      -- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006C9") =>
      -- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006CA") =>
      -- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006CB") =>
      -- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006CC") =>
      -- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006CD") =>
      -- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006CE") =>
      -- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006CF") =>
      -- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006D0") =>
      -- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006D1") =>
      -- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006D2") =>
      -- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006D3") =>
      -- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006D4") =>
      -- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006D5") =>
      -- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006D6") =>
      -- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006D7") =>
      -- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006D8") =>
      -- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006D9") =>
      -- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006DA") =>
      -- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006DB") =>
      -- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006DC") =>
      -- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006DD") =>
      -- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006DE") =>
      -- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006DF") =>
      -- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006E0") =>
      -- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006E1") =>
      -- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006E2") =>
      -- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006E3") =>
      -- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006E4") =>
      -- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006E5") =>
      -- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006E6") =>
      -- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006E7") =>
      -- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006E8") =>
      -- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006E9") =>
      -- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006EA") =>
      -- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006EB") =>
      -- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006EC") =>
      -- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006ED") =>
      -- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006EE") =>
      -- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006EF") =>
      -- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006F0") =>
      -- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006F1") =>
      -- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006F2") =>
      -- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006F3") =>
      -- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006F4") =>
      -- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006F5") =>
      -- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006F6") =>
      -- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006F7") =>
      -- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006F8") =>
      -- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006F9") =>
      -- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006FA") =>
      -- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006FB") =>
      -- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000006FC") =>
      -- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000006FD") =>
      -- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000006FE") =>
      -- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000006FF") =>
      -- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000700") =>
      -- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000701") =>
      -- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000702") =>
      -- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000703") =>
      -- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000704") =>
      -- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000705") =>
      -- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000706") =>
      -- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000707") =>
      -- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000708") =>
      -- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000709") =>
      -- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000070A") =>
      -- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000070B") =>
      -- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000070C") =>
      -- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000070D") =>
      -- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000070E") =>
      -- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000070F") =>
      -- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000710") =>
      -- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000711") =>
      -- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000712") =>
      -- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000713") =>
      -- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000714") =>
      -- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000715") =>
      -- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000716") =>
      -- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000717") =>
      -- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000718") =>
      -- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000719") =>
      -- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000071A") =>
      -- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000071B") =>
      -- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000071C") =>
      -- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000071D") =>
      -- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000071E") =>
      -- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000071F") =>
      -- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000720") =>
      -- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000721") =>
      -- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000722") =>
      -- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000723") =>
      -- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000724") =>
      -- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000725") =>
      -- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000726") =>
      -- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000727") =>
      -- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000728") =>
      -- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000729") =>
      -- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000072A") =>
      -- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000072B") =>
      -- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000072C") =>
      -- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000072D") =>
      -- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000072E") =>
      -- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000072F") =>
      -- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000730") =>
      -- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000731") =>
      -- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000732") =>
      -- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000733") =>
      -- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000734") =>
      -- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000735") =>
      -- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000736") =>
      -- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000737") =>
      -- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000738") =>
      -- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000739") =>
      -- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000073A") =>
      -- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000073B") =>
      -- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000073C") =>
      -- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000073D") =>
      -- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000073E") =>
      -- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000073F") =>
      -- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000740") =>
      -- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000741") =>
      -- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000742") =>
      -- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000743") =>
      -- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000744") =>
      -- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000745") =>
      -- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000746") =>
      -- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000747") =>
      -- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000748") =>
      -- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000749") =>
      -- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000074A") =>
      -- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000074B") =>
      -- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000074C") =>
      -- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000074D") =>
      -- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000074E") =>
      -- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000074F") =>
      -- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000750") =>
      -- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000751") =>
      -- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000752") =>
      -- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000753") =>
      -- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000754") =>
      -- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000755") =>
      -- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000756") =>
      -- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000757") =>
      -- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000758") =>
      -- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000759") =>
      -- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000075A") =>
      -- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000075B") =>
      -- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000075C") =>
      -- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000075D") =>
      -- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000075E") =>
      -- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000075F") =>
      -- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000760") =>
      -- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000761") =>
      -- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000762") =>
      -- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000763") =>
      -- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000764") =>
      -- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000765") =>
      -- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000766") =>
      -- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000767") =>
      -- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000768") =>
      -- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000769") =>
      -- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000076A") =>
      -- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000076B") =>
      -- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000076C") =>
      -- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000076D") =>
      -- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000076E") =>
      -- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000076F") =>
      -- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000770") =>
      -- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000771") =>
      -- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000772") =>
      -- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000773") =>
      -- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000774") =>
      -- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000775") =>
      -- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000776") =>
      -- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000777") =>
      -- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000778") =>
      -- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000779") =>
      -- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000077A") =>
      -- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000077B") =>
      -- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000077C") =>
      -- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000077D") =>
      -- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000077E") =>
      -- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000077F") =>
      -- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000780") =>
      -- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000781") =>
      -- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000782") =>
      -- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000783") =>
      -- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000784") =>
      -- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000785") =>
      -- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000786") =>
      -- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000787") =>
      -- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000788") =>
      -- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000789") =>
      -- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000078A") =>
      -- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000078B") =>
      -- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000078C") =>
      -- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000078D") =>
      -- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000078E") =>
      -- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000078F") =>
      -- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000790") =>
      -- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000791") =>
      -- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000792") =>
      -- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000793") =>
      -- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000794") =>
      -- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000795") =>
      -- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000796") =>
      -- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000797") =>
      -- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000798") =>
      -- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000799") =>
      -- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000079A") =>
      -- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000079B") =>
      -- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000079C") =>
      -- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000079D") =>
      -- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000079E") =>
      -- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000079F") =>
      -- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007A0") =>
      -- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007A1") =>
      -- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007A2") =>
      -- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007A3") =>
      -- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007A4") =>
      -- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007A5") =>
      -- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007A6") =>
      -- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007A7") =>
      -- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007A8") =>
      -- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007A9") =>
      -- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007AA") =>
      -- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007AB") =>
      -- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007AC") =>
      -- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007AD") =>
      -- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007AE") =>
      -- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007AF") =>
      -- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007B0") =>
      -- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007B1") =>
      -- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007B2") =>
      -- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007B3") =>
      -- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007B4") =>
      -- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007B5") =>
      -- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007B6") =>
      -- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007B7") =>
      -- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007B8") =>
      -- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007B9") =>
      -- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007BA") =>
      -- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007BB") =>
      -- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007BC") =>
      -- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007BD") =>
      -- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007BE") =>
      -- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007BF") =>
      -- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007C0") =>
      -- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007C1") =>
      -- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007C2") =>
      -- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007C3") =>
      -- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007C4") =>
      -- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007C5") =>
      -- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007C6") =>
      -- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007C7") =>
      -- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007C8") =>
      -- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007C9") =>
      -- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007CA") =>
      -- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007CB") =>
      -- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007CC") =>
      -- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007CD") =>
      -- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007CE") =>
      -- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007CF") =>
      -- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007D0") =>
      -- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007D1") =>
      -- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007D2") =>
      -- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007D3") =>
      -- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007D4") =>
      -- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007D5") =>
      -- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007D6") =>
      -- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007D7") =>
      -- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007D8") =>
      -- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007D9") =>
      -- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007DA") =>
      -- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007DB") =>
      -- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007DC") =>
      -- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007DD") =>
      -- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007DE") =>
      -- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007DF") =>
      -- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007E0") =>
      -- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007E1") =>
      -- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007E2") =>
      -- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007E3") =>
      -- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007E4") =>
      -- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007E5") =>
      -- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007E6") =>
      -- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007E7") =>
      -- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007E8") =>
      -- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007E9") =>
      -- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007EA") =>
      -- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007EB") =>
      -- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007EC") =>
      -- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007ED") =>
      -- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007EE") =>
      -- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007EF") =>
      -- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007F0") =>
      -- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007F1") =>
      -- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007F2") =>
      -- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007F3") =>
      -- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007F4") =>
      -- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007F5") =>
      -- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007F6") =>
      -- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007F7") =>
      -- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007F8") =>
      -- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007F9") =>
      -- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007FA") =>
      -- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007FB") =>
      -- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000007FC") =>
      -- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000007FD") =>
      -- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000007FE") =>
      -- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000007FF") =>
      -- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000800") =>
      -- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000801") =>
      -- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000802") =>
      -- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000803") =>
      -- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000804") =>
      -- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000805") =>
      -- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000806") =>
      -- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000807") =>
      -- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000808") =>
      -- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000809") =>
      -- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000080A") =>
      -- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000080B") =>
      -- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000080C") =>
      -- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000080D") =>
      -- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000080E") =>
      -- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000080F") =>
      -- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000810") =>
      -- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000811") =>
      -- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000812") =>
      -- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000813") =>
      -- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000814") =>
      -- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000815") =>
      -- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000816") =>
      -- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000817") =>
      -- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000818") =>
      -- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000819") =>
      -- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000081A") =>
      -- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000081B") =>
      -- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000081C") =>
      -- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000081D") =>
      -- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000081E") =>
      -- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000081F") =>
      -- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000820") =>
      -- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000821") =>
      -- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000822") =>
      -- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000823") =>
      -- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000824") =>
      -- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000825") =>
      -- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000826") =>
      -- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000827") =>
      -- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000828") =>
      -- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000829") =>
      -- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000082A") =>
      -- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000082B") =>
      -- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000082C") =>
      -- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000082D") =>
      -- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000082E") =>
      -- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000082F") =>
      -- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000830") =>
      -- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000831") =>
      -- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000832") =>
      -- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000833") =>
      -- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000834") =>
      -- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000835") =>
      -- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000836") =>
      -- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000837") =>
      -- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000838") =>
      -- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000839") =>
      -- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000083A") =>
      -- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000083B") =>
      -- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000083C") =>
      -- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000083D") =>
      -- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000083E") =>
      -- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000083F") =>
      -- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000840") =>
      -- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000841") =>
      -- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000842") =>
      -- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000843") =>
      -- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000844") =>
      -- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000845") =>
      -- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000846") =>
      -- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000847") =>
      -- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000848") =>
      -- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000849") =>
      -- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000084A") =>
      -- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000084B") =>
      -- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000084C") =>
      -- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000084D") =>
      -- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000084E") =>
      -- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000084F") =>
      -- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000850") =>
      -- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000851") =>
      -- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000852") =>
      -- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000853") =>
      -- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000854") =>
      -- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000855") =>
      -- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000856") =>
      -- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000857") =>
      -- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000858") =>
      -- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000859") =>
      -- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000085A") =>
      -- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000085B") =>
      -- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000085C") =>
      -- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000085D") =>
      -- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000085E") =>
      -- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000085F") =>
      -- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000860") =>
      -- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000861") =>
      -- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000862") =>
      -- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000863") =>
      -- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000864") =>
      -- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000865") =>
      -- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000866") =>
      -- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000867") =>
      -- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000868") =>
      -- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000869") =>
      -- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000086A") =>
      -- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000086B") =>
      -- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000086C") =>
      -- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000086D") =>
      -- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000086E") =>
      -- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000086F") =>
      -- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000870") =>
      -- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000871") =>
      -- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000872") =>
      -- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000873") =>
      -- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000874") =>
      -- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000875") =>
      -- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000876") =>
      -- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000877") =>
      -- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000878") =>
      -- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000879") =>
      -- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000087A") =>
      -- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000087B") =>
      -- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000087C") =>
      -- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000087D") =>
      -- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000087E") =>
      -- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000087F") =>
      -- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000880") =>
      -- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000881") =>
      -- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000882") =>
      -- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000883") =>
      -- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000884") =>
      -- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000885") =>
      -- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000886") =>
      -- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000887") =>
      -- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000888") =>
      -- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000889") =>
      -- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000088A") =>
      -- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000088B") =>
      -- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000088C") =>
      -- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000088D") =>
      -- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000088E") =>
      -- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000088F") =>
      -- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000890") =>
      -- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000891") =>
      -- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000892") =>
      -- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000893") =>
      -- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000894") =>
      -- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000895") =>
      -- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000896") =>
      -- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000897") =>
      -- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000898") =>
      -- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000899") =>
      -- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000089A") =>
      -- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000089B") =>
      -- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000089C") =>
      -- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000089D") =>
      -- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000089E") =>
      -- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000089F") =>
      -- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008A0") =>
      -- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008A1") =>
      -- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008A2") =>
      -- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008A3") =>
      -- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008A4") =>
      -- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008A5") =>
      -- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008A6") =>
      -- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008A7") =>
      -- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008A8") =>
      -- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008A9") =>
      -- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008AA") =>
      -- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008AB") =>
      -- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008AC") =>
      -- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008AD") =>
      -- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008AE") =>
      -- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008AF") =>
      -- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008B0") =>
      -- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008B1") =>
      -- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008B2") =>
      -- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008B3") =>
      -- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008B4") =>
      -- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008B5") =>
      -- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008B6") =>
      -- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008B7") =>
      -- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008B8") =>
      -- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008B9") =>
      -- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008BA") =>
      -- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008BB") =>
      -- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008BC") =>
      -- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008BD") =>
      -- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008BE") =>
      -- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008BF") =>
      -- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008C0") =>
      -- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008C1") =>
      -- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008C2") =>
      -- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008C3") =>
      -- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008C4") =>
      -- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008C5") =>
      -- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008C6") =>
      -- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008C7") =>
      -- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008C8") =>
      -- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008C9") =>
      -- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008CA") =>
      -- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008CB") =>
      -- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008CC") =>
      -- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008CD") =>
      -- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008CE") =>
      -- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008CF") =>
      -- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008D0") =>
      -- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008D1") =>
      -- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008D2") =>
      -- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008D3") =>
      -- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008D4") =>
      -- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008D5") =>
      -- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008D6") =>
      -- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008D7") =>
      -- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008D8") =>
      -- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008D9") =>
      -- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008DA") =>
      -- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008DB") =>
      -- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008DC") =>
      -- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008DD") =>
      -- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008DE") =>
      -- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008DF") =>
      -- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008E0") =>
      -- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008E1") =>
      -- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008E2") =>
      -- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008E3") =>
      -- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008E4") =>
      -- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008E5") =>
      -- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008E6") =>
      -- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008E7") =>
      -- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008E8") =>
      -- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008E9") =>
      -- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008EA") =>
      -- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008EB") =>
      -- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008EC") =>
      -- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008ED") =>
      -- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008EE") =>
      -- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008EF") =>
      -- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008F0") =>
      -- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008F1") =>
      -- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008F2") =>
      -- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008F3") =>
      -- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008F4") =>
      -- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008F5") =>
      -- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008F6") =>
      -- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008F7") =>
      -- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008F8") =>
      -- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008F9") =>
      -- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008FA") =>
      -- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008FB") =>
      -- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000008FC") =>
      -- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000008FD") =>
      -- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000008FE") =>
      -- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000008FF") =>
      -- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000900") =>
      -- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000901") =>
      -- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000902") =>
      -- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000903") =>
      -- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000904") =>
      -- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000905") =>
      -- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000906") =>
      -- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000907") =>
      -- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000908") =>
      -- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000909") =>
      -- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000090A") =>
      -- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000090B") =>
      -- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000090C") =>
      -- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000090D") =>
      -- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000090E") =>
      -- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000090F") =>
      -- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000910") =>
      -- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000911") =>
      -- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000912") =>
      -- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000913") =>
      -- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000914") =>
      -- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000915") =>
      -- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000916") =>
      -- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000917") =>
      -- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000918") =>
      -- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000919") =>
      -- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000091A") =>
      -- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000091B") =>
      -- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000091C") =>
      -- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000091D") =>
      -- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000091E") =>
      -- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000091F") =>
      -- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000920") =>
      -- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000921") =>
      -- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000922") =>
      -- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000923") =>
      -- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000924") =>
      -- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000925") =>
      -- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000926") =>
      -- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000927") =>
      -- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000928") =>
      -- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000929") =>
      -- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000092A") =>
      -- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000092B") =>
      -- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000092C") =>
      -- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000092D") =>
      -- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000092E") =>
      -- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000092F") =>
      -- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000930") =>
      -- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000931") =>
      -- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000932") =>
      -- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000933") =>
      -- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000934") =>
      -- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000935") =>
      -- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000936") =>
      -- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000937") =>
      -- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000938") =>
      -- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000939") =>
      -- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000093A") =>
      -- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000093B") =>
      -- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000093C") =>
      -- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000093D") =>
      -- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000093E") =>
      -- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000093F") =>
      -- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000940") =>
      -- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000941") =>
      -- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000942") =>
      -- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000943") =>
      -- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000944") =>
      -- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000945") =>
      -- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000946") =>
      -- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000947") =>
      -- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000948") =>
      -- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000949") =>
      -- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000094A") =>
      -- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000094B") =>
      -- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000094C") =>
      -- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000094D") =>
      -- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000094E") =>
      -- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000094F") =>
      -- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000950") =>
      -- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000951") =>
      -- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000952") =>
      -- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000953") =>
      -- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000954") =>
      -- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000955") =>
      -- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000956") =>
      -- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000957") =>
      -- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000958") =>
      -- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000959") =>
      -- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000095A") =>
      -- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000095B") =>
      -- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000095C") =>
      -- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000095D") =>
      -- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000095E") =>
      -- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000095F") =>
      -- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000960") =>
      -- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000961") =>
      -- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000962") =>
      -- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000963") =>
      -- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000964") =>
      -- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000965") =>
      -- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000966") =>
      -- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000967") =>
      -- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000968") =>
      -- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000969") =>
      -- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000096A") =>
      -- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000096B") =>
      -- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000096C") =>
      -- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000096D") =>
      -- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000096E") =>
      -- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000096F") =>
      -- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000970") =>
      -- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000971") =>
      -- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000972") =>
      -- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000973") =>
      -- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000974") =>
      -- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000975") =>
      -- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000976") =>
      -- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000977") =>
      -- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000978") =>
      -- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000979") =>
      -- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000097A") =>
      -- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000097B") =>
      -- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000097C") =>
      -- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000097D") =>
      -- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000097E") =>
      -- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000097F") =>
      -- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000980") =>
      -- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000981") =>
      -- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000982") =>
      -- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000983") =>
      -- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000984") =>
      -- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000985") =>
      -- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000986") =>
      -- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000987") =>
      -- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000988") =>
      -- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000989") =>
      -- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000098A") =>
      -- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000098B") =>
      -- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000098C") =>
      -- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000098D") =>
      -- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000098E") =>
      -- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000098F") =>
      -- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000990") =>
      -- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000991") =>
      -- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000992") =>
      -- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000993") =>
      -- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000994") =>
      -- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000995") =>
      -- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000996") =>
      -- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000997") =>
      -- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000998") =>
      -- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000999") =>
      -- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000099A") =>
      -- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000099B") =>
      -- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"0000099C") =>
      -- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"0000099D") =>
      -- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"0000099E") =>
      -- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"0000099F") =>
      -- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009A0") =>
      -- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009A1") =>
      -- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009A2") =>
      -- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009A3") =>
      -- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009A4") =>
      -- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009A5") =>
      -- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009A6") =>
      -- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009A7") =>
      -- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009A8") =>
      -- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009A9") =>
      -- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009AA") =>
      -- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009AB") =>
      -- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009AC") =>
      -- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009AD") =>
      -- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009AE") =>
      -- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009AF") =>
      -- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009B0") =>
      -- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009B1") =>
      -- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009B2") =>
      -- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009B3") =>
      -- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009B4") =>
      -- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009B5") =>
      -- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009B6") =>
      -- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009B7") =>
      -- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009B8") =>
      -- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009B9") =>
      -- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009BA") =>
      -- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009BB") =>
      -- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009BC") =>
      -- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009BD") =>
      -- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009BE") =>
      -- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009BF") =>
      -- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009C0") =>
      -- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009C1") =>
      -- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009C2") =>
      -- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009C3") =>
      -- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009C4") =>
      -- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009C5") =>
      -- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009C6") =>
      -- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009C7") =>
      -- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009C8") =>
      -- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009C9") =>
      -- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009CA") =>
      -- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009CB") =>
      -- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009CC") =>
      -- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009CD") =>
      -- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009CE") =>
      -- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009CF") =>
      -- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009D0") =>
      -- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009D1") =>
      -- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009D2") =>
      -- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009D3") =>
      -- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009D4") =>
      -- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009D5") =>
      -- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009D6") =>
      -- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009D7") =>
      -- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009D8") =>
      -- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009D9") =>
      -- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009DA") =>
      -- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009DB") =>
      -- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009DC") =>
      -- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009DD") =>
      -- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009DE") =>
      -- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009DF") =>
      -- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009E0") =>
      -- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009E1") =>
      -- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009E2") =>
      -- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009E3") =>
      -- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009E4") =>
      -- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009E5") =>
      -- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009E6") =>
      -- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009E7") =>
      -- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009E8") =>
      -- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009E9") =>
      -- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009EA") =>
      -- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009EB") =>
      -- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009EC") =>
      -- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009ED") =>
      -- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009EE") =>
      -- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009EF") =>
      -- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009F0") =>
      -- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009F1") =>
      -- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009F2") =>
      -- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009F3") =>
      -- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009F4") =>
      -- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009F5") =>
      -- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009F6") =>
      -- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009F7") =>
      -- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009F8") =>
      -- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009F9") =>
      -- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009FA") =>
      -- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009FB") =>
      -- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"000009FC") =>
      -- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"000009FD") =>
      -- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"000009FE") =>
      -- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"000009FF") =>
      -- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A00") =>
      -- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A01") =>
      -- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A02") =>
      -- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A03") =>
      -- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A04") =>
      -- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A05") =>
      -- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A06") =>
      -- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A07") =>
      -- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A08") =>
      -- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A09") =>
      -- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A0A") =>
      -- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A0B") =>
      -- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A0C") =>
      -- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A0D") =>
      -- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A0E") =>
      -- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A0F") =>
      -- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A10") =>
      -- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A11") =>
      -- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A12") =>
      -- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A13") =>
      -- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A14") =>
      -- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A15") =>
      -- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A16") =>
      -- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A17") =>
      -- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A18") =>
      -- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A19") =>
      -- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A1A") =>
      -- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A1B") =>
      -- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A1C") =>
      -- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A1D") =>
      -- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A1E") =>
      -- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A1F") =>
      -- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A20") =>
      -- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A21") =>
      -- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A22") =>
      -- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A23") =>
      -- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A24") =>
      -- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A25") =>
      -- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A26") =>
      -- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A27") =>
      -- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A28") =>
      -- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A29") =>
      -- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A2A") =>
      -- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A2B") =>
      -- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A2C") =>
      -- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A2D") =>
      -- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A2E") =>
      -- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A2F") =>
      -- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A30") =>
      -- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A31") =>
      -- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A32") =>
      -- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A33") =>
      -- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A34") =>
      -- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A35") =>
      -- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A36") =>
      -- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A37") =>
      -- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A38") =>
      -- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A39") =>
      -- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A3A") =>
      -- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A3B") =>
      -- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A3C") =>
      -- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A3D") =>
      -- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A3E") =>
      -- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A3F") =>
      -- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A40") =>
      -- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A41") =>
      -- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A42") =>
      -- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A43") =>
      -- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A44") =>
      -- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A45") =>
      -- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A46") =>
      -- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A47") =>
      -- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A48") =>
      -- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A49") =>
      -- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A4A") =>
      -- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A4B") =>
      -- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A4C") =>
      -- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A4D") =>
      -- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A4E") =>
      -- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A4F") =>
      -- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A50") =>
      -- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A51") =>
      -- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A52") =>
      -- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A53") =>
      -- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A54") =>
      -- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A55") =>
      -- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A56") =>
      -- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A57") =>
      -- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A58") =>
      -- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A59") =>
      -- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A5A") =>
      -- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A5B") =>
      -- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A5C") =>
      -- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A5D") =>
      -- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A5E") =>
      -- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A5F") =>
      -- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A60") =>
      -- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A61") =>
      -- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A62") =>
      -- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A63") =>
      -- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A64") =>
      -- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A65") =>
      -- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A66") =>
      -- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A67") =>
      -- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A68") =>
      -- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A69") =>
      -- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A6A") =>
      -- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A6B") =>
      -- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A6C") =>
      -- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A6D") =>
      -- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A6E") =>
      -- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A6F") =>
      -- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A70") =>
      -- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A71") =>
      -- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A72") =>
      -- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A73") =>
      -- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A74") =>
      -- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A75") =>
      -- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A76") =>
      -- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A77") =>
      -- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A78") =>
      -- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A79") =>
      -- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A7A") =>
      -- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A7B") =>
      -- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A7C") =>
      -- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A7D") =>
      -- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A7E") =>
      -- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A7F") =>
      -- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A80") =>
      -- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A81") =>
      -- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A82") =>
      -- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A83") =>
      -- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A84") =>
      -- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A85") =>
      -- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A86") =>
      -- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A87") =>
      -- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A88") =>
      -- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A89") =>
      -- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A8A") =>
      -- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A8B") =>
      -- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A8C") =>
      -- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A8D") =>
      -- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A8E") =>
      -- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A8F") =>
      -- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A90") =>
      -- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A91") =>
      -- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A92") =>
      -- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A93") =>
      -- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A94") =>
      -- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A95") =>
      -- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A96") =>
      -- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A97") =>
      -- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A98") =>
      -- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A99") =>
      -- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A9A") =>
      -- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A9B") =>
      -- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000A9C") =>
      -- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000A9D") =>
      -- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000A9E") =>
      -- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000A9F") =>
      -- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AA0") =>
      -- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AA1") =>
      -- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AA2") =>
      -- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AA3") =>
      -- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AA4") =>
      -- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AA5") =>
      -- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AA6") =>
      -- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AA7") =>
      -- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AA8") =>
      -- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AA9") =>
      -- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AAA") =>
      -- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AAB") =>
      -- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AAC") =>
      -- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AAD") =>
      -- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AAE") =>
      -- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AAF") =>
      -- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AB0") =>
      -- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AB1") =>
      -- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AB2") =>
      -- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AB3") =>
      -- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AB4") =>
      -- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AB5") =>
      -- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AB6") =>
      -- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AB7") =>
      -- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AB8") =>
      -- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AB9") =>
      -- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ABA") =>
      -- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ABB") =>
      -- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ABC") =>
      -- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ABD") =>
      -- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ABE") =>
      -- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ABF") =>
      -- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AC0") =>
      -- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AC1") =>
      -- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AC2") =>
      -- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AC3") =>
      -- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AC4") =>
      -- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AC5") =>
      -- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AC6") =>
      -- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AC7") =>
      -- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AC8") =>
      -- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AC9") =>
      -- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ACA") =>
      -- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ACB") =>
      -- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ACC") =>
      -- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ACD") =>
      -- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ACE") =>
      -- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ACF") =>
      -- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AD0") =>
      -- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AD1") =>
      -- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AD2") =>
      -- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AD3") =>
      -- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AD4") =>
      -- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AD5") =>
      -- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AD6") =>
      -- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AD7") =>
      -- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AD8") =>
      -- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AD9") =>
      -- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ADA") =>
      -- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ADB") =>
      -- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ADC") =>
      -- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ADD") =>
      -- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ADE") =>
      -- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ADF") =>
      -- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AE0") =>
      -- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AE1") =>
      -- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AE2") =>
      -- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AE3") =>
      -- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AE4") =>
      -- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AE5") =>
      -- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AE6") =>
      -- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AE7") =>
      -- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AE8") =>
      -- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AE9") =>
      -- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AEA") =>
      -- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AEB") =>
      -- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AEC") =>
      -- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AED") =>
      -- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AEE") =>
      -- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AEF") =>
      -- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AF0") =>
      -- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AF1") =>
      -- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AF2") =>
      -- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AF3") =>
      -- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AF4") =>
      -- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AF5") =>
      -- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AF6") =>
      -- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AF7") =>
      -- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AF8") =>
      -- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AF9") =>
      -- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AFA") =>
      -- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AFB") =>
      -- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000AFC") =>
      -- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000AFD") =>
      -- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000AFE") =>
      -- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000AFF") =>
      -- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B00") =>
      -- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B01") =>
      -- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B02") =>
      -- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B03") =>
      -- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B04") =>
      -- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B05") =>
      -- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B06") =>
      -- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B07") =>
      -- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B08") =>
      -- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B09") =>
      -- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B0A") =>
      -- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B0B") =>
      -- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B0C") =>
      -- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B0D") =>
      -- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B0E") =>
      -- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B0F") =>
      -- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B10") =>
      -- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B11") =>
      -- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B12") =>
      -- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B13") =>
      -- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B14") =>
      -- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B15") =>
      -- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B16") =>
      -- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B17") =>
      -- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B18") =>
      -- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B19") =>
      -- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B1A") =>
      -- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B1B") =>
      -- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B1C") =>
      -- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B1D") =>
      -- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B1E") =>
      -- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B1F") =>
      -- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B20") =>
      -- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B21") =>
      -- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B22") =>
      -- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B23") =>
      -- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B24") =>
      -- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B25") =>
      -- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B26") =>
      -- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B27") =>
      -- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B28") =>
      -- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B29") =>
      -- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B2A") =>
      -- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B2B") =>
      -- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B2C") =>
      -- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B2D") =>
      -- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B2E") =>
      -- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B2F") =>
      -- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B30") =>
      -- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B31") =>
      -- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B32") =>
      -- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B33") =>
      -- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B34") =>
      -- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B35") =>
      -- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B36") =>
      -- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B37") =>
      -- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B38") =>
      -- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B39") =>
      -- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B3A") =>
      -- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B3B") =>
      -- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B3C") =>
      -- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B3D") =>
      -- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B3E") =>
      -- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B3F") =>
      -- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B40") =>
      -- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B41") =>
      -- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B42") =>
      -- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B43") =>
      -- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B44") =>
      -- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B45") =>
      -- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B46") =>
      -- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B47") =>
      -- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B48") =>
      -- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B49") =>
      -- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B4A") =>
      -- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B4B") =>
      -- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B4C") =>
      -- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B4D") =>
      -- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B4E") =>
      -- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B4F") =>
      -- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B50") =>
      -- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B51") =>
      -- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B52") =>
      -- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B53") =>
      -- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B54") =>
      -- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B55") =>
      -- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B56") =>
      -- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B57") =>
      -- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B58") =>
      -- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B59") =>
      -- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B5A") =>
      -- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B5B") =>
      -- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B5C") =>
      -- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B5D") =>
      -- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B5E") =>
      -- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B5F") =>
      -- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B60") =>
      -- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B61") =>
      -- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B62") =>
      -- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B63") =>
      -- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B64") =>
      -- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B65") =>
      -- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B66") =>
      -- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B67") =>
      -- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B68") =>
      -- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B69") =>
      -- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B6A") =>
      -- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B6B") =>
      -- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B6C") =>
      -- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B6D") =>
      -- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B6E") =>
      -- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B6F") =>
      -- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B70") =>
      -- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B71") =>
      -- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B72") =>
      -- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B73") =>
      -- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B74") =>
      -- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B75") =>
      -- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B76") =>
      -- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B77") =>
      -- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B78") =>
      -- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B79") =>
      -- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B7A") =>
      -- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B7B") =>
      -- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B7C") =>
      -- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B7D") =>
      -- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B7E") =>
      -- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B7F") =>
      -- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B80") =>
      -- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B81") =>
      -- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B82") =>
      -- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B83") =>
      -- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B84") =>
      -- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B85") =>
      -- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B86") =>
      -- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B87") =>
      -- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B88") =>
      -- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B89") =>
      -- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B8A") =>
      -- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B8B") =>
      -- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B8C") =>
      -- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B8D") =>
      -- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B8E") =>
      -- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B8F") =>
      -- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B90") =>
      -- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B91") =>
      -- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B92") =>
      -- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B93") =>
      -- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B94") =>
      -- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B95") =>
      -- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B96") =>
      -- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B97") =>
      -- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B98") =>
      -- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B99") =>
      -- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B9A") =>
      -- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B9B") =>
      -- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000B9C") =>
      -- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000B9D") =>
      -- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000B9E") =>
      -- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000B9F") =>
      -- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BA0") =>
      -- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BA1") =>
      -- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BA2") =>
      -- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BA3") =>
      -- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BA4") =>
      -- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BA5") =>
      -- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BA6") =>
      -- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BA7") =>
      -- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BA8") =>
      -- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BA9") =>
      -- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BAA") =>
      -- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BAB") =>
      -- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BAC") =>
      -- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BAD") =>
      -- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BAE") =>
      -- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BAF") =>
      -- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BB0") =>
      -- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BB1") =>
      -- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BB2") =>
      -- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BB3") =>
      -- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BB4") =>
      -- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BB5") =>
      -- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BB6") =>
      -- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BB7") =>
      -- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BB8") =>
      -- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BB9") =>
      -- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BBA") =>
      -- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BBB") =>
      -- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BBC") =>
      -- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BBD") =>
      -- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BBE") =>
      -- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BBF") =>
      -- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BC0") =>
      -- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BC1") =>
      -- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BC2") =>
      -- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BC3") =>
      -- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BC4") =>
      -- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BC5") =>
      -- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BC6") =>
      -- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BC7") =>
      -- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BC8") =>
      -- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BC9") =>
      -- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BCA") =>
      -- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BCB") =>
      -- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BCC") =>
      -- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BCD") =>
      -- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BCE") =>
      -- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BCF") =>
      -- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BD0") =>
      -- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BD1") =>
      -- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BD2") =>
      -- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BD3") =>
      -- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BD4") =>
      -- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BD5") =>
      -- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BD6") =>
      -- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BD7") =>
      -- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BD8") =>
      -- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BD9") =>
      -- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BDA") =>
      -- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BDB") =>
      -- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BDC") =>
      -- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BDD") =>
      -- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BDE") =>
      -- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BDF") =>
      -- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BE0") =>
      -- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BE1") =>
      -- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BE2") =>
      -- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BE3") =>
      -- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BE4") =>
      -- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BE5") =>
      -- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BE6") =>
      -- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BE7") =>
      -- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BE8") =>
      -- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BE9") =>
      -- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BEA") =>
      -- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BEB") =>
      -- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BEC") =>
      -- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BED") =>
      -- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BEE") =>
      -- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BEF") =>
      -- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BF0") =>
      -- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BF1") =>
      -- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BF2") =>
      -- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BF3") =>
      -- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BF4") =>
      -- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BF5") =>
      -- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BF6") =>
      -- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BF7") =>
      -- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BF8") =>
      -- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BF9") =>
      -- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BFA") =>
      -- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BFB") =>
      -- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000BFC") =>
      -- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000BFD") =>
      -- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000BFE") =>
      -- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000BFF") =>
      -- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C00") =>
      -- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C01") =>
      -- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C02") =>
      -- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C03") =>
      -- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C04") =>
      -- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C05") =>
      -- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C06") =>
      -- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C07") =>
      -- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C08") =>
      -- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C09") =>
      -- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C0A") =>
      -- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C0B") =>
      -- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C0C") =>
      -- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C0D") =>
      -- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C0E") =>
      -- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C0F") =>
      -- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C10") =>
      -- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C11") =>
      -- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C12") =>
      -- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C13") =>
      -- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C14") =>
      -- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C15") =>
      -- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C16") =>
      -- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C17") =>
      -- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C18") =>
      -- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C19") =>
      -- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C1A") =>
      -- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C1B") =>
      -- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C1C") =>
      -- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C1D") =>
      -- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C1E") =>
      -- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C1F") =>
      -- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C20") =>
      -- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C21") =>
      -- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C22") =>
      -- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C23") =>
      -- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C24") =>
      -- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C25") =>
      -- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C26") =>
      -- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C27") =>
      -- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C28") =>
      -- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C29") =>
      -- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C2A") =>
      -- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C2B") =>
      -- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C2C") =>
      -- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C2D") =>
      -- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C2E") =>
      -- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C2F") =>
      -- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C30") =>
      -- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C31") =>
      -- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C32") =>
      -- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C33") =>
      -- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C34") =>
      -- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C35") =>
      -- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C36") =>
      -- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C37") =>
      -- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C38") =>
      -- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C39") =>
      -- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C3A") =>
      -- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C3B") =>
      -- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C3C") =>
      -- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C3D") =>
      -- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C3E") =>
      -- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C3F") =>
      -- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C40") =>
      -- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C41") =>
      -- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C42") =>
      -- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C43") =>
      -- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C44") =>
      -- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C45") =>
      -- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C46") =>
      -- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C47") =>
      -- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C48") =>
      -- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C49") =>
      -- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C4A") =>
      -- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C4B") =>
      -- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C4C") =>
      -- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C4D") =>
      -- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C4E") =>
      -- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C4F") =>
      -- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C50") =>
      -- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C51") =>
      -- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C52") =>
      -- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C53") =>
      -- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C54") =>
      -- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C55") =>
      -- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C56") =>
      -- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C57") =>
      -- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C58") =>
      -- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C59") =>
      -- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C5A") =>
      -- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C5B") =>
      -- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C5C") =>
      -- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C5D") =>
      -- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C5E") =>
      -- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C5F") =>
      -- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C60") =>
      -- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C61") =>
      -- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C62") =>
      -- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C63") =>
      -- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C64") =>
      -- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C65") =>
      -- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C66") =>
      -- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C67") =>
      -- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C68") =>
      -- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C69") =>
      -- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C6A") =>
      -- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C6B") =>
      -- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C6C") =>
      -- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C6D") =>
      -- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C6E") =>
      -- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C6F") =>
      -- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C70") =>
      -- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C71") =>
      -- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C72") =>
      -- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C73") =>
      -- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C74") =>
      -- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C75") =>
      -- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C76") =>
      -- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C77") =>
      -- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C78") =>
      -- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C79") =>
      -- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C7A") =>
      -- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C7B") =>
      -- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C7C") =>
      -- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C7D") =>
      -- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C7E") =>
      -- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C7F") =>
      -- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C80") =>
      -- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C81") =>
      -- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C82") =>
      -- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C83") =>
      -- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C84") =>
      -- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C85") =>
      -- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C86") =>
      -- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C87") =>
      -- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C88") =>
      -- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C89") =>
      -- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C8A") =>
      -- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C8B") =>
      -- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C8C") =>
      -- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C8D") =>
      -- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C8E") =>
      -- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C8F") =>
      -- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C90") =>
      -- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C91") =>
      -- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C92") =>
      -- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C93") =>
      -- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C94") =>
      -- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C95") =>
      -- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C96") =>
      -- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C97") =>
      -- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C98") =>
      -- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C99") =>
      -- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C9A") =>
      -- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C9B") =>
      -- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000C9C") =>
      -- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000C9D") =>
      -- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000C9E") =>
      -- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000C9F") =>
      -- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CA0") =>
      -- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CA1") =>
      -- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CA2") =>
      -- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CA3") =>
      -- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CA4") =>
      -- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CA5") =>
      -- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CA6") =>
      -- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CA7") =>
      -- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CA8") =>
      -- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CA9") =>
      -- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CAA") =>
      -- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CAB") =>
      -- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CAC") =>
      -- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CAD") =>
      -- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CAE") =>
      -- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CAF") =>
      -- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CB0") =>
      -- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CB1") =>
      -- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CB2") =>
      -- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CB3") =>
      -- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CB4") =>
      -- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CB5") =>
      -- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CB6") =>
      -- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CB7") =>
      -- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CB8") =>
      -- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CB9") =>
      -- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CBA") =>
      -- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CBB") =>
      -- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CBC") =>
      -- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CBD") =>
      -- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CBE") =>
      -- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CBF") =>
      -- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CC0") =>
      -- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CC1") =>
      -- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CC2") =>
      -- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CC3") =>
      -- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CC4") =>
      -- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CC5") =>
      -- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CC6") =>
      -- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CC7") =>
      -- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CC8") =>
      -- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CC9") =>
      -- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CCA") =>
      -- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CCB") =>
      -- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CCC") =>
      -- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CCD") =>
      -- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CCE") =>
      -- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CCF") =>
      -- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CD0") =>
      -- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CD1") =>
      -- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CD2") =>
      -- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CD3") =>
      -- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CD4") =>
      -- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CD5") =>
      -- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CD6") =>
      -- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CD7") =>
      -- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CD8") =>
      -- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CD9") =>
      -- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CDA") =>
      -- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CDB") =>
      -- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CDC") =>
      -- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CDD") =>
      -- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CDE") =>
      -- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CDF") =>
      -- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CE0") =>
      -- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CE1") =>
      -- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CE2") =>
      -- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CE3") =>
      -- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CE4") =>
      -- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CE5") =>
      -- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CE6") =>
      -- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CE7") =>
      -- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CE8") =>
      -- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CE9") =>
      -- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CEA") =>
      -- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CEB") =>
      -- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CEC") =>
      -- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CED") =>
      -- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CEE") =>
      -- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CEF") =>
      -- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CF0") =>
      -- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CF1") =>
      -- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CF2") =>
      -- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CF3") =>
      -- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CF4") =>
      -- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CF5") =>
      -- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CF6") =>
      -- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CF7") =>
      -- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CF8") =>
      -- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CF9") =>
      -- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CFA") =>
      -- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CFB") =>
      -- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000CFC") =>
      -- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000CFD") =>
      -- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000CFE") =>
      -- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000CFF") =>
      -- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D00") =>
      -- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D01") =>
      -- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D02") =>
      -- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D03") =>
      -- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D04") =>
      -- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D05") =>
      -- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D06") =>
      -- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D07") =>
      -- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D08") =>
      -- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D09") =>
      -- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D0A") =>
      -- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D0B") =>
      -- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D0C") =>
      -- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D0D") =>
      -- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D0E") =>
      -- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D0F") =>
      -- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D10") =>
      -- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D11") =>
      -- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D12") =>
      -- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D13") =>
      -- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D14") =>
      -- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D15") =>
      -- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D16") =>
      -- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D17") =>
      -- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D18") =>
      -- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D19") =>
      -- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D1A") =>
      -- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D1B") =>
      -- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D1C") =>
      -- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D1D") =>
      -- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D1E") =>
      -- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D1F") =>
      -- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D20") =>
      -- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D21") =>
      -- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D22") =>
      -- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D23") =>
      -- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D24") =>
      -- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D25") =>
      -- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D26") =>
      -- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D27") =>
      -- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D28") =>
      -- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D29") =>
      -- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D2A") =>
      -- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D2B") =>
      -- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D2C") =>
      -- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D2D") =>
      -- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D2E") =>
      -- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D2F") =>
      -- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D30") =>
      -- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D31") =>
      -- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D32") =>
      -- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D33") =>
      -- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D34") =>
      -- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D35") =>
      -- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D36") =>
      -- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D37") =>
      -- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D38") =>
      -- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D39") =>
      -- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D3A") =>
      -- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D3B") =>
      -- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D3C") =>
      -- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D3D") =>
      -- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D3E") =>
      -- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D3F") =>
      -- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D40") =>
      -- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D41") =>
      -- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D42") =>
      -- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D43") =>
      -- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D44") =>
      -- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D45") =>
      -- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D46") =>
      -- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D47") =>
      -- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D48") =>
      -- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D49") =>
      -- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D4A") =>
      -- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D4B") =>
      -- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D4C") =>
      -- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D4D") =>
      -- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D4E") =>
      -- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D4F") =>
      -- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D50") =>
      -- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D51") =>
      -- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D52") =>
      -- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D53") =>
      -- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D54") =>
      -- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D55") =>
      -- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D56") =>
      -- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D57") =>
      -- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D58") =>
      -- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D59") =>
      -- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D5A") =>
      -- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D5B") =>
      -- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D5C") =>
      -- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D5D") =>
      -- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D5E") =>
      -- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D5F") =>
      -- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D60") =>
      -- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D61") =>
      -- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D62") =>
      -- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D63") =>
      -- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D64") =>
      -- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D65") =>
      -- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D66") =>
      -- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D67") =>
      -- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D68") =>
      -- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D69") =>
      -- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D6A") =>
      -- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D6B") =>
      -- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D6C") =>
      -- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D6D") =>
      -- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D6E") =>
      -- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D6F") =>
      -- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D70") =>
      -- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D71") =>
      -- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D72") =>
      -- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D73") =>
      -- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D74") =>
      -- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D75") =>
      -- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D76") =>
      -- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D77") =>
      -- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D78") =>
      -- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D79") =>
      -- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D7A") =>
      -- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D7B") =>
      -- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D7C") =>
      -- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D7D") =>
      -- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D7E") =>
      -- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D7F") =>
      -- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D80") =>
      -- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D81") =>
      -- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D82") =>
      -- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D83") =>
      -- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D84") =>
      -- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D85") =>
      -- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D86") =>
      -- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D87") =>
      -- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D88") =>
      -- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D89") =>
      -- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D8A") =>
      -- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D8B") =>
      -- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D8C") =>
      -- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D8D") =>
      -- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D8E") =>
      -- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D8F") =>
      -- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D90") =>
      -- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D91") =>
      -- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D92") =>
      -- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D93") =>
      -- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D94") =>
      -- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D95") =>
      -- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D96") =>
      -- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D97") =>
      -- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D98") =>
      -- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D99") =>
      -- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D9A") =>
      -- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D9B") =>
      -- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000D9C") =>
      -- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000D9D") =>
      -- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000D9E") =>
      -- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000D9F") =>
      -- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DA0") =>
      -- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DA1") =>
      -- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DA2") =>
      -- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DA3") =>
      -- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DA4") =>
      -- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DA5") =>
      -- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DA6") =>
      -- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DA7") =>
      -- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DA8") =>
      -- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DA9") =>
      -- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DAA") =>
      -- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DAB") =>
      -- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DAC") =>
      -- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DAD") =>
      -- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DAE") =>
      -- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DAF") =>
      -- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DB0") =>
      -- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DB1") =>
      -- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DB2") =>
      -- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DB3") =>
      -- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DB4") =>
      -- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DB5") =>
      -- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DB6") =>
      -- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DB7") =>
      -- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DB8") =>
      -- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DB9") =>
      -- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DBA") =>
      -- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DBB") =>
      -- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DBC") =>
      -- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DBD") =>
      -- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DBE") =>
      -- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DBF") =>
      -- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DC0") =>
      -- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DC1") =>
      -- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DC2") =>
      -- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DC3") =>
      -- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DC4") =>
      -- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DC5") =>
      -- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DC6") =>
      -- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DC7") =>
      -- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DC8") =>
      -- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DC9") =>
      -- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DCA") =>
      -- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DCB") =>
      -- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DCC") =>
      -- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DCD") =>
      -- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DCE") =>
      -- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DCF") =>
      -- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DD0") =>
      -- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DD1") =>
      -- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DD2") =>
      -- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DD3") =>
      -- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DD4") =>
      -- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DD5") =>
      -- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DD6") =>
      -- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DD7") =>
      -- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DD8") =>
      -- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DD9") =>
      -- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DDA") =>
      -- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DDB") =>
      -- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DDC") =>
      -- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DDD") =>
      -- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DDE") =>
      -- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DDF") =>
      -- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DE0") =>
      -- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DE1") =>
      -- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DE2") =>
      -- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DE3") =>
      -- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DE4") =>
      -- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DE5") =>
      -- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DE6") =>
      -- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DE7") =>
      -- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DE8") =>
      -- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DE9") =>
      -- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DEA") =>
      -- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DEB") =>
      -- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DEC") =>
      -- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DED") =>
      -- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DEE") =>
      -- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DEF") =>
      -- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DF0") =>
      -- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DF1") =>
      -- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DF2") =>
      -- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DF3") =>
      -- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DF4") =>
      -- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DF5") =>
      -- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DF6") =>
      -- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DF7") =>
      -- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DF8") =>
      -- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DF9") =>
      -- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DFA") =>
      -- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DFB") =>
      -- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000DFC") =>
      -- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000DFD") =>
      -- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000DFE") =>
      -- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000DFF") =>
      -- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E00") =>
      -- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E01") =>
      -- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E02") =>
      -- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E03") =>
      -- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E04") =>
      -- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E05") =>
      -- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E06") =>
      -- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E07") =>
      -- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E08") =>
      -- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E09") =>
      -- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E0A") =>
      -- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E0B") =>
      -- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E0C") =>
      -- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E0D") =>
      -- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E0E") =>
      -- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E0F") =>
      -- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E10") =>
      -- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E11") =>
      -- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E12") =>
      -- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E13") =>
      -- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E14") =>
      -- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E15") =>
      -- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E16") =>
      -- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E17") =>
      -- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E18") =>
      -- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E19") =>
      -- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E1A") =>
      -- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E1B") =>
      -- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E1C") =>
      -- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E1D") =>
      -- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E1E") =>
      -- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E1F") =>
      -- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E20") =>
      -- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E21") =>
      -- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E22") =>
      -- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E23") =>
      -- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E24") =>
      -- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E25") =>
      -- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E26") =>
      -- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E27") =>
      -- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E28") =>
      -- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E29") =>
      -- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E2A") =>
      -- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E2B") =>
      -- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E2C") =>
      -- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E2D") =>
      -- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E2E") =>
      -- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E2F") =>
      -- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E30") =>
      -- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E31") =>
      -- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E32") =>
      -- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E33") =>
      -- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E34") =>
      -- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E35") =>
      -- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E36") =>
      -- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E37") =>
      -- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E38") =>
      -- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E39") =>
      -- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E3A") =>
      -- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E3B") =>
      -- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E3C") =>
      -- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E3D") =>
      -- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E3E") =>
      -- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E3F") =>
      -- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E40") =>
      -- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E41") =>
      -- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E42") =>
      -- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E43") =>
      -- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E44") =>
      -- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E45") =>
      -- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E46") =>
      -- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E47") =>
      -- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E48") =>
      -- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E49") =>
      -- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E4A") =>
      -- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E4B") =>
      -- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E4C") =>
      -- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E4D") =>
      -- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E4E") =>
      -- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E4F") =>
      -- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E50") =>
      -- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E51") =>
      -- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E52") =>
      -- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E53") =>
      -- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E54") =>
      -- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E55") =>
      -- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E56") =>
      -- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E57") =>
      -- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E58") =>
      -- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E59") =>
      -- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E5A") =>
      -- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E5B") =>
      -- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E5C") =>
      -- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E5D") =>
      -- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E5E") =>
      -- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E5F") =>
      -- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E60") =>
      -- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E61") =>
      -- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E62") =>
      -- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E63") =>
      -- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E64") =>
      -- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E65") =>
      -- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E66") =>
      -- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E67") =>
      -- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E68") =>
      -- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E69") =>
      -- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E6A") =>
      -- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E6B") =>
      -- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E6C") =>
      -- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E6D") =>
      -- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E6E") =>
      -- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E6F") =>
      -- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E70") =>
      -- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E71") =>
      -- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E72") =>
      -- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E73") =>
      -- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E74") =>
      -- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E75") =>
      -- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E76") =>
      -- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E77") =>
      -- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E78") =>
      -- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E79") =>
      -- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E7A") =>
      -- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E7B") =>
      -- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E7C") =>
      -- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E7D") =>
      -- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E7E") =>
      -- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E7F") =>
      -- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E80") =>
      -- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E81") =>
      -- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E82") =>
      -- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E83") =>
      -- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E84") =>
      -- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E85") =>
      -- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E86") =>
      -- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E87") =>
      -- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E88") =>
      -- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E89") =>
      -- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E8A") =>
      -- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E8B") =>
      -- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E8C") =>
      -- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E8D") =>
      -- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E8E") =>
      -- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E8F") =>
      -- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E90") =>
      -- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E91") =>
      -- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E92") =>
      -- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E93") =>
      -- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E94") =>
      -- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E95") =>
      -- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E96") =>
      -- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E97") =>
      -- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E98") =>
      -- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E99") =>
      -- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E9A") =>
      -- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E9B") =>
      -- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000E9C") =>
      -- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000E9D") =>
      -- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000E9E") =>
      -- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000E9F") =>
      -- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EA0") =>
      -- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EA1") =>
      -- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EA2") =>
      -- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EA3") =>
      -- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EA4") =>
      -- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EA5") =>
      -- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EA6") =>
      -- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EA7") =>
      -- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EA8") =>
      -- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EA9") =>
      -- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EAA") =>
      -- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EAB") =>
      -- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EAC") =>
      -- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EAD") =>
      -- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EAE") =>
      -- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EAF") =>
      -- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EB0") =>
      -- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EB1") =>
      -- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EB2") =>
      -- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EB3") =>
      -- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EB4") =>
      -- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EB5") =>
      -- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EB6") =>
      -- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EB7") =>
      -- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EB8") =>
      -- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EB9") =>
      -- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EBA") =>
      -- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EBB") =>
      -- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EBC") =>
      -- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EBD") =>
      -- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EBE") =>
      -- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EBF") =>
      -- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EC0") =>
      -- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EC1") =>
      -- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EC2") =>
      -- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EC3") =>
      -- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EC4") =>
      -- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EC5") =>
      -- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EC6") =>
      -- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EC7") =>
      -- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EC8") =>
      -- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EC9") =>
      -- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ECA") =>
      -- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ECB") =>
      -- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ECC") =>
      -- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ECD") =>
      -- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ECE") =>
      -- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ECF") =>
      -- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ED0") =>
      -- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ED1") =>
      -- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ED2") =>
      -- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ED3") =>
      -- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ED4") =>
      -- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ED5") =>
      -- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000ED6") =>
      -- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000ED7") =>
      -- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000ED8") =>
      -- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000ED9") =>
      -- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EDA") =>
      -- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EDB") =>
      -- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EDC") =>
      -- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EDD") =>
      -- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EDE") =>
      -- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EDF") =>
      -- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EE0") =>
      -- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EE1") =>
      -- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EE2") =>
      -- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EE3") =>
      -- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EE4") =>
      -- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EE5") =>
      -- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EE6") =>
      -- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EE7") =>
      -- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EE8") =>
      -- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EE9") =>
      -- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EEA") =>
      -- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EEB") =>
      -- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EEC") =>
      -- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EED") =>
      -- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EEE") =>
      -- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EEF") =>
      -- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EF0") =>
      -- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EF1") =>
      -- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EF2") =>
      -- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EF3") =>
      -- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EF4") =>
      -- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EF5") =>
      -- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EF6") =>
      -- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EF7") =>
      -- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EF8") =>
      -- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EF9") =>
      -- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EFA") =>
      -- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EFB") =>
      -- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000EFC") =>
      -- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000EFD") =>
      -- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000EFE") =>
      -- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000EFF") =>
      -- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F00") =>
      -- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F01") =>
      -- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F02") =>
      -- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F03") =>
      -- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F04") =>
      -- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F05") =>
      -- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F06") =>
      -- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F07") =>
      -- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F08") =>
      -- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F09") =>
      -- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F0A") =>
      -- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F0B") =>
      -- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F0C") =>
      -- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F0D") =>
      -- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F0E") =>
      -- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F0F") =>
      -- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F10") =>
      -- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F11") =>
      -- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F12") =>
      -- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F13") =>
      -- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F14") =>
      -- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F15") =>
      -- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F16") =>
      -- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F17") =>
      -- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F18") =>
      -- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F19") =>
      -- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F1A") =>
      -- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F1B") =>
      -- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F1C") =>
      -- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F1D") =>
      -- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F1E") =>
      -- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F1F") =>
      -- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F20") =>
      -- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F21") =>
      -- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F22") =>
      -- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F23") =>
      -- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F24") =>
      -- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F25") =>
      -- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F26") =>
      -- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F27") =>
      -- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F28") =>
      -- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F29") =>
      -- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F2A") =>
      -- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F2B") =>
      -- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F2C") =>
      -- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F2D") =>
      -- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F2E") =>
      -- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F2F") =>
      -- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F30") =>
      -- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F31") =>
      -- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F32") =>
      -- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F33") =>
      -- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F34") =>
      -- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F35") =>
      -- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F36") =>
      -- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F37") =>
      -- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F38") =>
      -- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F39") =>
      -- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F3A") =>
      -- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F3B") =>
      -- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F3C") =>
      -- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F3D") =>
      -- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F3E") =>
      -- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F3F") =>
      -- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F40") =>
      -- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F41") =>
      -- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F42") =>
      -- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F43") =>
      -- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F44") =>
      -- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F45") =>
      -- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F46") =>
      -- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F47") =>
      -- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F48") =>
      -- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F49") =>
      -- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F4A") =>
      -- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F4B") =>
      -- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F4C") =>
      -- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F4D") =>
      -- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F4E") =>
      -- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F4F") =>
      -- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F50") =>
      -- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F51") =>
      -- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F52") =>
      -- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F53") =>
      -- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F54") =>
      -- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F55") =>
      -- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F56") =>
      -- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F57") =>
      -- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F58") =>
      -- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F59") =>
      -- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F5A") =>
      -- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F5B") =>
      -- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F5C") =>
      -- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F5D") =>
      -- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F5E") =>
      -- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F5F") =>
      -- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F60") =>
      -- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F61") =>
      -- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F62") =>
      -- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F63") =>
      -- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F64") =>
      -- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F65") =>
      -- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F66") =>
      -- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F67") =>
      -- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F68") =>
      -- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F69") =>
      -- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F6A") =>
      -- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F6B") =>
      -- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F6C") =>
      -- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F6D") =>
      -- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F6E") =>
      -- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F6F") =>
      -- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F70") =>
      -- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F71") =>
      -- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F72") =>
      -- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F73") =>
      -- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F74") =>
      -- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F75") =>
      -- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F76") =>
      -- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F77") =>
      -- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F78") =>
      -- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F79") =>
      -- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F7A") =>
      -- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F7B") =>
      -- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F7C") =>
      -- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F7D") =>
      -- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F7E") =>
      -- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F7F") =>
      -- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F80") =>
      -- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F81") =>
      -- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F82") =>
      -- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F83") =>
      -- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F84") =>
      -- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F85") =>
      -- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F86") =>
      -- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F87") =>
      -- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F88") =>
      -- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F89") =>
      -- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F8A") =>
      -- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F8B") =>
      -- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F8C") =>
      -- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F8D") =>
      -- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F8E") =>
      -- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F8F") =>
      -- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F90") =>
      -- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F91") =>
      -- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F92") =>
      -- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F93") =>
      -- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F94") =>
      -- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F95") =>
      -- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F96") =>
      -- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F97") =>
      -- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F98") =>
      -- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F99") =>
      -- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F9A") =>
      -- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F9B") =>
      -- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000F9C") =>
      -- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000F9D") =>
      -- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000F9E") =>
      -- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000F9F") =>
      -- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FA0") =>
      -- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FA1") =>
      -- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FA2") =>
      -- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FA3") =>
      -- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FA4") =>
      -- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FA5") =>
      -- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FA6") =>
      -- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FA7") =>
      -- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FA8") =>
      -- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FA9") =>
      -- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FAA") =>
      -- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FAB") =>
      -- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FAC") =>
      -- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FAD") =>
      -- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FAE") =>
      -- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FAF") =>
      -- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FB0") =>
      -- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FB1") =>
      -- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FB2") =>
      -- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FB3") =>
      -- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FB4") =>
      -- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FB5") =>
      -- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FB6") =>
      -- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FB7") =>
      -- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FB8") =>
      -- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FB9") =>
      -- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FBA") =>
      -- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FBB") =>
      -- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FBC") =>
      -- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FBD") =>
      -- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FBE") =>
      -- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FBF") =>
      -- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FC0") =>
      -- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FC1") =>
      -- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FC2") =>
      -- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FC3") =>
      -- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FC4") =>
      -- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FC5") =>
      -- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FC6") =>
      -- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FC7") =>
      -- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FC8") =>
      -- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FC9") =>
      -- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FCA") =>
      -- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FCB") =>
      -- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FCC") =>
      -- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FCD") =>
      -- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FCE") =>
      -- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FCF") =>
      -- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FD0") =>
      -- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FD1") =>
      -- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FD2") =>
      -- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FD3") =>
      -- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FD4") =>
      -- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FD5") =>
      -- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FD6") =>
      -- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FD7") =>
      -- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FD8") =>
      -- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FD9") =>
      -- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FDA") =>
      -- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FDB") =>
      -- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FDC") =>
      -- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FDD") =>
      -- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FDE") =>
      -- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FDF") =>
      -- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FE0") =>
      -- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FE1") =>
      -- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FE2") =>
      -- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FE3") =>
      -- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FE4") =>
      -- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FE5") =>
      -- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FE6") =>
      -- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FE7") =>
      -- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FE8") =>
      -- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FE9") =>
      -- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FEA") =>
      -- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FEB") =>
      -- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FEC") =>
      -- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FED") =>
      -- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FEE") =>
      -- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FEF") =>
      -- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FF0") =>
      -- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FF1") =>
      -- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FF2") =>
      -- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FF3") =>
      -- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FF4") =>
      -- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FF5") =>
      -- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FF6") =>
      -- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FF7") =>
      -- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FF8") =>
      -- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FF9") =>
      -- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FFA") =>
      -- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FFB") =>
      -- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when (x"00000FFC") =>
      -- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(31 downto 24) <= fee_rmap_i.writedata;

  when (x"00000FFD") =>
      -- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(23 downto 16) <= fee_rmap_i.writedata;

  when (x"00000FFE") =>
      -- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(15 downto 8) <= fee_rmap_i.writedata;

  when (x"00000FFF") =>
      -- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(7 downto 0) <= fee_rmap_i.writedata;

  when others =>
    null;

end case;

		end procedure p_ffee_aeb_mem_wr;

		-- p_avalon_mm_rmap_write

		procedure p_avs_writedata(write_address_i : t_farm_avalon_mm_rmap_ffee_aeb_address) is
		begin

-- Registers Write Data
case (write_address_i) is
  -- Case for access to all registers address

  when (16#000#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;

  when (16#001#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "NEW_STATE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.new_state <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;

  when (16#002#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "SET_STATE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.set_state <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#003#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "AEB_RESET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.aeb_reset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#004#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_1 <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;

  when (16#005#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_DATA_RD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_data_rd <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#006#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_WR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_wr <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#007#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "ADC_CFG_RD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.adc_cfg_rd <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#008#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "DAC_WR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.dac_wr <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#009#) =>
      -- AEB Critical Configuration Area Register "AEB_CONTROL" : "RESERVED_2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_2(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_control.reserved_2(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_0 <= avalon_mm_rmap_i.writedata(21 downto 16);
    end if;

  when (16#00A#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "WATCH-DOG_DIS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.watchdog_dis <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#00B#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "INT_SYNC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.int_sync <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#00C#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_1 <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#00D#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP_CDS_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp_cds_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#00E#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP2_CAL_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp2_cal_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#00F#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "VASP1_CAL_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.vasp1_cal_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#010#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG" : "RESERVED_2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_2(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config.reserved_2(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#011#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_KEY" : "KEY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_key.key(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#012#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_SW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_sw <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#013#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;

  when (16#014#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#015#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#016#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VAN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_van1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#017#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCLK" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vclk <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#018#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "SW_VCCD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.sw_vccd <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#019#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_VASP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_vasp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01A#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01B#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_PIX_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_pix_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01C#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_PIX_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_pix_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01D#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_ADC_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_adc_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01E#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_ADC_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_adc_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#01F#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP2_RESET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp2_reset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#020#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "VASP1_RESET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.vasp1_reset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#021#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "OVERRIDE_ADC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.override_adc <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#022#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_EN_P5V0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_en_p5v0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#023#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_EN_P5V0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_en_p5v0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#024#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "PT1000_CAL_ON_N" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.pt1000_cal_on_n <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#025#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "EN_V_MUX_N" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.en_v_mux_n <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#026#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC2_PWDN_N" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc2_pwdn_n <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#027#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC1_PWDN_N" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc1_pwdn_n <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#028#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "ADC_CLK_EN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.adc_clk_en <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#029#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_AIT" : "RESERVED_2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_ait.reserved_2 <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_CCDID" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_ccdid <= avalon_mm_rmap_i.writedata(9 downto 8);
    end if;
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_COLS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_cols(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_cols(13 downto 8) <= avalon_mm_rmap_i.writedata(29 downto 24);
    end if;

  when (16#02A#) =>
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.reserved <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "AEB_CONFIG_PATTERN" : "PATTERN_ROWS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_rows(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_aeb_config_pattern.pattern_rows(13 downto 8) <= avalon_mm_rmap_i.writedata(29 downto 24);
    end if;

  when (16#02B#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP_CFG_ADDR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp_cfg_addr <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_CFG_DATA" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_cfg_data <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_CFG_DATA" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_cfg_data <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.reserved <= avalon_mm_rmap_i.writedata(26 downto 24);
    end if;

  when (16#02C#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP2_SELECT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp2_select <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#02D#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "VASP1_SELECT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.vasp1_select <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#02E#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "CALIBRATION_START" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.calibration_start <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#02F#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_READ_START" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_read_start <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#030#) =>
      -- AEB Critical Configuration Area Register "VASP_I2C_CONTROL" : "I2C_WRITE_START" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_vasp_i2c_control.i2c_write_start <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#031#) =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_0 <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VOG" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vog(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vog(11 downto 8) <= avalon_mm_rmap_i.writedata(27 downto 24);
    end if;

  when (16#032#) =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.reserved_1 <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "DAC_CONFIG_1" : "DAC_VRD" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vrd(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_1.dac_vrd(11 downto 8) <= avalon_mm_rmap_i.writedata(27 downto 24);
    end if;

  when (16#033#) =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_0 <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "DAC_VOD" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.dac_vod(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.dac_vod(11 downto 8) <= avalon_mm_rmap_i.writedata(27 downto 24);
    end if;

  when (16#034#) =>
      -- AEB Critical Configuration Area Register "DAC_CONFIG_2" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_1(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_dac_config_2.reserved_1(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#035#) =>
      -- AEB Critical Configuration Area Register "RESERVED_20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#036#) =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCCD_ON" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vccd_on <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VCLK_ON" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_vclk_on <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN1_ON" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van1_on <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG1" : "TIME_VAN2_ON" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config1.time_van2_on <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#037#) =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN3_ON" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van3_on <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCCD_OFF" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vccd_off <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VCLK_OFF" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_vclk_off <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG2" : "TIME_VAN1_OFF" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config2.time_van1_off <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#038#) =>
      -- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN2_OFF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van2_off <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Critical Configuration Area Register "PWR_CONFIG3" : "TIME_VAN3_OFF" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_pwr_config3.time_van3_off <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#039#) =>
      -- AEB Critical Configuration Area Register "RESERVED_30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03A#) =>
      -- AEB Critical Configuration Area Register "RESERVED_34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03B#) =>
      -- AEB Critical Configuration Area Register "RESERVED_38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03C#) =>
      -- AEB Critical Configuration Area Register "RESERVED_3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03D#) =>
      -- AEB Critical Configuration Area Register "RESERVED_40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03E#) =>
      -- AEB Critical Configuration Area Register "RESERVED_44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#03F#) =>
      -- AEB Critical Configuration Area Register "RESERVED_48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#040#) =>
      -- AEB Critical Configuration Area Register "RESERVED_4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#041#) =>
      -- AEB Critical Configuration Area Register "RESERVED_50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#042#) =>
      -- AEB Critical Configuration Area Register "RESERVED_54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#043#) =>
      -- AEB Critical Configuration Area Register "RESERVED_58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#044#) =>
      -- AEB Critical Configuration Area Register "RESERVED_5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#045#) =>
      -- AEB Critical Configuration Area Register "RESERVED_60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#046#) =>
      -- AEB Critical Configuration Area Register "RESERVED_64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#047#) =>
      -- AEB Critical Configuration Area Register "RESERVED_68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#048#) =>
      -- AEB Critical Configuration Area Register "RESERVED_6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#049#) =>
      -- AEB Critical Configuration Area Register "RESERVED_70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04A#) =>
      -- AEB Critical Configuration Area Register "RESERVED_74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04B#) =>
      -- AEB Critical Configuration Area Register "RESERVED_78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04C#) =>
      -- AEB Critical Configuration Area Register "RESERVED_7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04D#) =>
      -- AEB Critical Configuration Area Register "RESERVED_80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04E#) =>
      -- AEB Critical Configuration Area Register "RESERVED_84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#04F#) =>
      -- AEB Critical Configuration Area Register "RESERVED_88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#050#) =>
      -- AEB Critical Configuration Area Register "RESERVED_8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#051#) =>
      -- AEB Critical Configuration Area Register "RESERVED_90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#052#) =>
      -- AEB Critical Configuration Area Register "RESERVED_94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#053#) =>
      -- AEB Critical Configuration Area Register "RESERVED_98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#054#) =>
      -- AEB Critical Configuration Area Register "RESERVED_9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#055#) =>
      -- AEB Critical Configuration Area Register "RESERVED_A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#056#) =>
      -- AEB Critical Configuration Area Register "RESERVED_A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#057#) =>
      -- AEB Critical Configuration Area Register "RESERVED_A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#058#) =>
      -- AEB Critical Configuration Area Register "RESERVED_AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#059#) =>
      -- AEB Critical Configuration Area Register "RESERVED_B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05A#) =>
      -- AEB Critical Configuration Area Register "RESERVED_B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05B#) =>
      -- AEB Critical Configuration Area Register "RESERVED_B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05C#) =>
      -- AEB Critical Configuration Area Register "RESERVED_BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05D#) =>
      -- AEB Critical Configuration Area Register "RESERVED_C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05E#) =>
      -- AEB Critical Configuration Area Register "RESERVED_C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#05F#) =>
      -- AEB Critical Configuration Area Register "RESERVED_C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#060#) =>
      -- AEB Critical Configuration Area Register "RESERVED_CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#061#) =>
      -- AEB Critical Configuration Area Register "RESERVED_D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#062#) =>
      -- AEB Critical Configuration Area Register "RESERVED_D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#063#) =>
      -- AEB Critical Configuration Area Register "RESERVED_D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#064#) =>
      -- AEB Critical Configuration Area Register "RESERVED_DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#065#) =>
      -- AEB Critical Configuration Area Register "RESERVED_E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#066#) =>
      -- AEB Critical Configuration Area Register "RESERVED_E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#067#) =>
      -- AEB Critical Configuration Area Register "RESERVED_E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#068#) =>
      -- AEB Critical Configuration Area Register "RESERVED_EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#069#) =>
      -- AEB Critical Configuration Area Register "RESERVED_F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#06A#) =>
      -- AEB Critical Configuration Area Register "RESERVED_F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#06B#) =>
      -- AEB Critical Configuration Area Register "RESERVED_F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#06C#) =>
      -- AEB Critical Configuration Area Register "RESERVED_FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_crit_cfg_reserved_fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#06D#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#06E#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SPIRST" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.spirst <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#06F#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "MUXMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.muxmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#070#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "BYPAS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.bypas <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#071#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CLKENB" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.clkenb <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#072#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "CHOP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.chop <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#073#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "STAT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.stat <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#074#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#075#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "IDLMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.idlmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#076#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.dly <= avalon_mm_rmap_i.writedata(2 downto 0);
    end if;
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "SBCS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.sbcs <= avalon_mm_rmap_i.writedata(9 downto 8);
    end if;
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DRATE" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.drate <= avalon_mm_rmap_i.writedata(17 downto 16);
    end if;
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINP" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainp <= avalon_mm_rmap_i.writedata(27 downto 24);
    end if;

  when (16#077#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "AINN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.ainn <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;
      -- AEB General Configuration Area Register "ADC1_CONFIG_1" : "DIFF" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_1.diff <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#078#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#079#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07A#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07B#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07C#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07D#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07E#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#07F#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#080#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN15" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain15 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#081#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN14" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain14 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#082#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN13" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain13 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#083#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN12" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain12 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#084#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN11" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain11 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#085#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN10" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain10 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#086#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN9" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain9 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#087#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "AIN8" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ain8 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#088#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;

  when (16#089#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "REF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.ref <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08A#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "GAIN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.gain <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08B#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "TEMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.temp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08C#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "VCC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.vcc <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08D#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08E#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "OFFSET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.offset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#08F#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#090#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#091#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#092#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#093#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#094#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#095#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#096#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_2" : "CIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_2.cio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#097#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#098#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#099#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09A#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09B#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09C#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09D#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09E#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "DIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.dio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#09F#) =>
      -- AEB General Configuration Area Register "ADC1_CONFIG_3" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc1_config_3.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#0A0#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A1#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SPIRST" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.spirst <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A2#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "MUXMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.muxmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A3#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "BYPAS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.bypas <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A4#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CLKENB" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.clkenb <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A5#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "CHOP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.chop <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A6#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "STAT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.stat <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A7#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A8#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "IDLMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.idlmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0A9#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.dly <= avalon_mm_rmap_i.writedata(2 downto 0);
    end if;
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "SBCS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.sbcs <= avalon_mm_rmap_i.writedata(9 downto 8);
    end if;
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DRATE" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.drate <= avalon_mm_rmap_i.writedata(17 downto 16);
    end if;
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINP" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainp <= avalon_mm_rmap_i.writedata(27 downto 24);
    end if;

  when (16#0AA#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "AINN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.ainn <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;
      -- AEB General Configuration Area Register "ADC2_CONFIG_1" : "DIFF" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_1.diff <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#0AB#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0AC#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0AD#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0AE#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0AF#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B0#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B1#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B2#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B3#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN15" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain15 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B4#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN14" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain14 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B5#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN13" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain13 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B6#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN12" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain12 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B7#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN11" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain11 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B8#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN10" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain10 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0B9#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN9" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain9 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0BA#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "AIN8" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ain8 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0BB#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;

  when (16#0BC#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "REF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.ref <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0BD#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "GAIN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.gain <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0BE#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "TEMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.temp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0BF#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "VCC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.vcc <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C0#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C1#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "OFFSET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.offset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C2#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C3#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C4#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C5#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C6#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C7#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C8#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0C9#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_2" : "CIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_2.cio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CA#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CB#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CC#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CD#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CE#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0CF#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D0#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D1#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "DIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.dio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D2#) =>
      -- AEB General Configuration Area Register "ADC2_CONFIG_3" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_adc2_config_3.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#0D3#) =>
      -- AEB General Configuration Area Register "RESERVED_118" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_118.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0D4#) =>
      -- AEB General Configuration Area Register "RESERVED_11C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_11c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0D5#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;

  when (16#0D6#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_CCD_ENABLE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ccd_enable <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D7#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPARE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_spare <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D8#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTLINE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstline <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0D9#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TSTFRM" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tstfrm <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DA#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_VASPCLAMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_vaspclamp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DB#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_PRECLAMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_preclamp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DC#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IG" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_ig <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DD#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_TG" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_tg <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DE#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_DG" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_dg <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0DF#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHIR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphir <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E0#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sw <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E1#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E2#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E3#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_RPHI1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_rphi1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E4#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E5#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E6#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E7#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_SPHI1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_sphi1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E8#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0E9#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0EA#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0EB#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "SEQ_OE_IPHI1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.seq_oe_iphi1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0EC#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0ED#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_1" : "ADC_CLK_DIV" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_1.adc_clk_div <= avalon_mm_rmap_i.writedata(6 downto 0);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_low_pos <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "ADC_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.adc_clk_high_pos <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_low_pos <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0EE#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_2" : "CDS_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_2.cds_clk_high_pos <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_low_pos <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHIR_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphir_clk_high_pos <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_low_pos <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0EF#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_3" : "RPHI1_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_3.rphi1_clk_high_pos <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_low_pos <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI2_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi2_clk_high_pos <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_low_pos <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0F0#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_4" : "RPHI3_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_4.rphi3_clk_high_pos <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_LOW_POS" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_low_pos <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "SW_CLK_HIGH_POS" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.sw_clk_high_pos <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#0F1#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_CTRL" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_ctrl <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0F2#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.reserved <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0F3#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_5" : "VASP_OUT_EN_POS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_en_pos(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_5.vasp_out_en_pos(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;

  when (16#0F4#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_CTRL_INV" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_ctrl_inv <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0F5#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0F6#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "VASP_OUT_DIS_POS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_dis_pos(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.vasp_out_dis_pos(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_6" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_1(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_6.reserved_1(15 downto 8) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0F7#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_7" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_7.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0F8#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#0F9#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_0 <= avalon_mm_rmap_i.writedata(1 downto 0);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "FT_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.ft_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.ft_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(29 downto 24);
    end if;

  when (16#0FA#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_ENABLED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_enabled <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0FB#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0FC#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_9" : "LT0_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_9.lt0_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;

  when (16#0FD#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_ENABLED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_enabled <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0FE#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#0FF#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT1_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt1_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;

  when (16#100#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_ENABLED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_enabled <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#101#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.reserved_1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#102#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_10" : "LT2_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_10.lt2_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;

  when (16#103#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_ENABLED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_enabled <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#104#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.reserved <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#105#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "LT3_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.lt3_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_11" : "PIX_LOOP_CNT_WORD_1" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.pix_loop_cnt_word_1(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_11.pix_loop_cnt_word_1(15 downto 8) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#106#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PIX_LOOP_CNT_WORD_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pix_loop_cnt_word_0(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pix_loop_cnt_word_0(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#107#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_ENABLED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_enabled <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#108#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.reserved <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#109#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_12" : "PC_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_12.pc_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_0 <= avalon_mm_rmap_i.writedata(17 downto 16);
    end if;

  when (16#10A#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT1_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int1_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int1_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.reserved_1 <= avalon_mm_rmap_i.writedata(17 downto 16);
    end if;

  when (16#10B#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_13" : "INT2_LOOP_CNT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int2_loop_cnt(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_13.int2_loop_cnt(13 downto 8) <= avalon_mm_rmap_i.writedata(13 downto 8);
    end if;
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_0" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_0 <= avalon_mm_rmap_i.writedata(22 downto 16);
    end if;

  when (16#10C#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "SPHI_INV" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.sphi_inv <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#10D#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_1 <= avalon_mm_rmap_i.writedata(6 downto 0);
    end if;

  when (16#10E#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RPHI_INV" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.rphi_inv <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#10F#) =>
      -- AEB General Configuration Area Register "SEQ_CONFIG_14" : "RESERVED_2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_2(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_seq_config_14.reserved_2(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;

  when (16#110#) =>
      -- AEB General Configuration Area Register "RESERVED_158" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_158.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#111#) =>
      -- AEB General Configuration Area Register "RESERVED_15C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_15c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#112#) =>
      -- AEB General Configuration Area Register "RESERVED_160" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_160.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#113#) =>
      -- AEB General Configuration Area Register "RESERVED_164" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_164.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#114#) =>
      -- AEB General Configuration Area Register "RESERVED_168" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_168.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#115#) =>
      -- AEB General Configuration Area Register "RESERVED_16C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_16c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#116#) =>
      -- AEB General Configuration Area Register "RESERVED_170" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_170.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#117#) =>
      -- AEB General Configuration Area Register "RESERVED_174" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_174.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#118#) =>
      -- AEB General Configuration Area Register "RESERVED_178" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_178.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#119#) =>
      -- AEB General Configuration Area Register "RESERVED_17C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_17c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11A#) =>
      -- AEB General Configuration Area Register "RESERVED_180" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_180.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11B#) =>
      -- AEB General Configuration Area Register "RESERVED_184" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_184.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11C#) =>
      -- AEB General Configuration Area Register "RESERVED_188" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_188.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11D#) =>
      -- AEB General Configuration Area Register "RESERVED_18C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_18c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11E#) =>
      -- AEB General Configuration Area Register "RESERVED_190" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_190.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#11F#) =>
      -- AEB General Configuration Area Register "RESERVED_194" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_194.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#120#) =>
      -- AEB General Configuration Area Register "RESERVED_198" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_198.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#121#) =>
      -- AEB General Configuration Area Register "RESERVED_19C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_19c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#122#) =>
      -- AEB General Configuration Area Register "RESERVED_1A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#123#) =>
      -- AEB General Configuration Area Register "RESERVED_1A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#124#) =>
      -- AEB General Configuration Area Register "RESERVED_1A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#125#) =>
      -- AEB General Configuration Area Register "RESERVED_1AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#126#) =>
      -- AEB General Configuration Area Register "RESERVED_1B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#127#) =>
      -- AEB General Configuration Area Register "RESERVED_1B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#128#) =>
      -- AEB General Configuration Area Register "RESERVED_1B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#129#) =>
      -- AEB General Configuration Area Register "RESERVED_1BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12A#) =>
      -- AEB General Configuration Area Register "RESERVED_1C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12B#) =>
      -- AEB General Configuration Area Register "RESERVED_1C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12C#) =>
      -- AEB General Configuration Area Register "RESERVED_1C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12D#) =>
      -- AEB General Configuration Area Register "RESERVED_1CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12E#) =>
      -- AEB General Configuration Area Register "RESERVED_1D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#12F#) =>
      -- AEB General Configuration Area Register "RESERVED_1D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#130#) =>
      -- AEB General Configuration Area Register "RESERVED_1D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#131#) =>
      -- AEB General Configuration Area Register "RESERVED_1DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#132#) =>
      -- AEB General Configuration Area Register "RESERVED_1E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#133#) =>
      -- AEB General Configuration Area Register "RESERVED_1E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#134#) =>
      -- AEB General Configuration Area Register "RESERVED_1E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#135#) =>
      -- AEB General Configuration Area Register "RESERVED_1EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#136#) =>
      -- AEB General Configuration Area Register "RESERVED_1F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#137#) =>
      -- AEB General Configuration Area Register "RESERVED_1F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#138#) =>
      -- AEB General Configuration Area Register "RESERVED_1F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#139#) =>
      -- AEB General Configuration Area Register "RESERVED_1FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_1fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13A#) =>
      -- AEB General Configuration Area Register "RESERVED_200" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_200.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13B#) =>
      -- AEB General Configuration Area Register "RESERVED_204" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_204.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13C#) =>
      -- AEB General Configuration Area Register "RESERVED_208" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_208.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13D#) =>
      -- AEB General Configuration Area Register "RESERVED_20C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_20c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13E#) =>
      -- AEB General Configuration Area Register "RESERVED_210" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_210.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#13F#) =>
      -- AEB General Configuration Area Register "RESERVED_214" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_214.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#140#) =>
      -- AEB General Configuration Area Register "RESERVED_218" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_218.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#141#) =>
      -- AEB General Configuration Area Register "RESERVED_21C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_21c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#142#) =>
      -- AEB General Configuration Area Register "RESERVED_220" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_220.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#143#) =>
      -- AEB General Configuration Area Register "RESERVED_224" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_224.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#144#) =>
      -- AEB General Configuration Area Register "RESERVED_228" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_228.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#145#) =>
      -- AEB General Configuration Area Register "RESERVED_22C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_22c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#146#) =>
      -- AEB General Configuration Area Register "RESERVED_230" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_230.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#147#) =>
      -- AEB General Configuration Area Register "RESERVED_234" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_234.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#148#) =>
      -- AEB General Configuration Area Register "RESERVED_238" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_238.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#149#) =>
      -- AEB General Configuration Area Register "RESERVED_23C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_23c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14A#) =>
      -- AEB General Configuration Area Register "RESERVED_240" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_240.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14B#) =>
      -- AEB General Configuration Area Register "RESERVED_244" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_244.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14C#) =>
      -- AEB General Configuration Area Register "RESERVED_248" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_248.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14D#) =>
      -- AEB General Configuration Area Register "RESERVED_24C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_24c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14E#) =>
      -- AEB General Configuration Area Register "RESERVED_250" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_250.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#14F#) =>
      -- AEB General Configuration Area Register "RESERVED_254" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_254.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#150#) =>
      -- AEB General Configuration Area Register "RESERVED_258" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_258.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#151#) =>
      -- AEB General Configuration Area Register "RESERVED_25C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_25c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#152#) =>
      -- AEB General Configuration Area Register "RESERVED_260" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_260.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#153#) =>
      -- AEB General Configuration Area Register "RESERVED_264" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_264.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#154#) =>
      -- AEB General Configuration Area Register "RESERVED_268" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_268.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#155#) =>
      -- AEB General Configuration Area Register "RESERVED_26C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_26c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#156#) =>
      -- AEB General Configuration Area Register "RESERVED_270" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_270.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#157#) =>
      -- AEB General Configuration Area Register "RESERVED_274" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_274.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#158#) =>
      -- AEB General Configuration Area Register "RESERVED_278" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_278.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#159#) =>
      -- AEB General Configuration Area Register "RESERVED_27C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_27c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15A#) =>
      -- AEB General Configuration Area Register "RESERVED_280" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_280.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15B#) =>
      -- AEB General Configuration Area Register "RESERVED_284" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_284.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15C#) =>
      -- AEB General Configuration Area Register "RESERVED_288" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_288.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15D#) =>
      -- AEB General Configuration Area Register "RESERVED_28C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_28c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15E#) =>
      -- AEB General Configuration Area Register "RESERVED_290" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_290.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#15F#) =>
      -- AEB General Configuration Area Register "RESERVED_294" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_294.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#160#) =>
      -- AEB General Configuration Area Register "RESERVED_298" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_298.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#161#) =>
      -- AEB General Configuration Area Register "RESERVED_29C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_29c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#162#) =>
      -- AEB General Configuration Area Register "RESERVED_2A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#163#) =>
      -- AEB General Configuration Area Register "RESERVED_2A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#164#) =>
      -- AEB General Configuration Area Register "RESERVED_2A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#165#) =>
      -- AEB General Configuration Area Register "RESERVED_2AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#166#) =>
      -- AEB General Configuration Area Register "RESERVED_2B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#167#) =>
      -- AEB General Configuration Area Register "RESERVED_2B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#168#) =>
      -- AEB General Configuration Area Register "RESERVED_2B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#169#) =>
      -- AEB General Configuration Area Register "RESERVED_2BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16A#) =>
      -- AEB General Configuration Area Register "RESERVED_2C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16B#) =>
      -- AEB General Configuration Area Register "RESERVED_2C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16C#) =>
      -- AEB General Configuration Area Register "RESERVED_2C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16D#) =>
      -- AEB General Configuration Area Register "RESERVED_2CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16E#) =>
      -- AEB General Configuration Area Register "RESERVED_2D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#16F#) =>
      -- AEB General Configuration Area Register "RESERVED_2D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#170#) =>
      -- AEB General Configuration Area Register "RESERVED_2D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#171#) =>
      -- AEB General Configuration Area Register "RESERVED_2DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#172#) =>
      -- AEB General Configuration Area Register "RESERVED_2E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#173#) =>
      -- AEB General Configuration Area Register "RESERVED_2E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#174#) =>
      -- AEB General Configuration Area Register "RESERVED_2E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#175#) =>
      -- AEB General Configuration Area Register "RESERVED_2EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#176#) =>
      -- AEB General Configuration Area Register "RESERVED_2F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#177#) =>
      -- AEB General Configuration Area Register "RESERVED_2F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#178#) =>
      -- AEB General Configuration Area Register "RESERVED_2F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#179#) =>
      -- AEB General Configuration Area Register "RESERVED_2FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_2fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17A#) =>
      -- AEB General Configuration Area Register "RESERVED_300" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_300.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17B#) =>
      -- AEB General Configuration Area Register "RESERVED_304" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_304.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17C#) =>
      -- AEB General Configuration Area Register "RESERVED_308" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_308.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17D#) =>
      -- AEB General Configuration Area Register "RESERVED_30C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_30c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17E#) =>
      -- AEB General Configuration Area Register "RESERVED_310" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_310.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#17F#) =>
      -- AEB General Configuration Area Register "RESERVED_314" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_314.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#180#) =>
      -- AEB General Configuration Area Register "RESERVED_318" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_318.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#181#) =>
      -- AEB General Configuration Area Register "RESERVED_31C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_31c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#182#) =>
      -- AEB General Configuration Area Register "RESERVED_320" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_320.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#183#) =>
      -- AEB General Configuration Area Register "RESERVED_324" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_324.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#184#) =>
      -- AEB General Configuration Area Register "RESERVED_328" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_328.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#185#) =>
      -- AEB General Configuration Area Register "RESERVED_32C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_32c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#186#) =>
      -- AEB General Configuration Area Register "RESERVED_330" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_330.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#187#) =>
      -- AEB General Configuration Area Register "RESERVED_334" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_334.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#188#) =>
      -- AEB General Configuration Area Register "RESERVED_338" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_338.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#189#) =>
      -- AEB General Configuration Area Register "RESERVED_33C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_33c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18A#) =>
      -- AEB General Configuration Area Register "RESERVED_340" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_340.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18B#) =>
      -- AEB General Configuration Area Register "RESERVED_344" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_344.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18C#) =>
      -- AEB General Configuration Area Register "RESERVED_348" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_348.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18D#) =>
      -- AEB General Configuration Area Register "RESERVED_34C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_34c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18E#) =>
      -- AEB General Configuration Area Register "RESERVED_350" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_350.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#18F#) =>
      -- AEB General Configuration Area Register "RESERVED_354" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_354.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#190#) =>
      -- AEB General Configuration Area Register "RESERVED_358" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_358.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#191#) =>
      -- AEB General Configuration Area Register "RESERVED_35C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_35c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#192#) =>
      -- AEB General Configuration Area Register "RESERVED_360" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_360.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#193#) =>
      -- AEB General Configuration Area Register "RESERVED_364" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_364.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#194#) =>
      -- AEB General Configuration Area Register "RESERVED_368" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_368.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#195#) =>
      -- AEB General Configuration Area Register "RESERVED_36C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_36c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#196#) =>
      -- AEB General Configuration Area Register "RESERVED_370" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_370.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#197#) =>
      -- AEB General Configuration Area Register "RESERVED_374" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_374.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#198#) =>
      -- AEB General Configuration Area Register "RESERVED_378" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_378.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#199#) =>
      -- AEB General Configuration Area Register "RESERVED_37C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_37c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19A#) =>
      -- AEB General Configuration Area Register "RESERVED_380" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_380.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19B#) =>
      -- AEB General Configuration Area Register "RESERVED_384" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_384.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19C#) =>
      -- AEB General Configuration Area Register "RESERVED_388" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_388.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19D#) =>
      -- AEB General Configuration Area Register "RESERVED_38C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_38c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19E#) =>
      -- AEB General Configuration Area Register "RESERVED_390" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_390.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#19F#) =>
      -- AEB General Configuration Area Register "RESERVED_394" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_394.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A0#) =>
      -- AEB General Configuration Area Register "RESERVED_398" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_398.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A1#) =>
      -- AEB General Configuration Area Register "RESERVED_39C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_39c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A2#) =>
      -- AEB General Configuration Area Register "RESERVED_3A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A3#) =>
      -- AEB General Configuration Area Register "RESERVED_3A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A4#) =>
      -- AEB General Configuration Area Register "RESERVED_3A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A5#) =>
      -- AEB General Configuration Area Register "RESERVED_3AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A6#) =>
      -- AEB General Configuration Area Register "RESERVED_3B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A7#) =>
      -- AEB General Configuration Area Register "RESERVED_3B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A8#) =>
      -- AEB General Configuration Area Register "RESERVED_3B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1A9#) =>
      -- AEB General Configuration Area Register "RESERVED_3BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AA#) =>
      -- AEB General Configuration Area Register "RESERVED_3C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AB#) =>
      -- AEB General Configuration Area Register "RESERVED_3C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AC#) =>
      -- AEB General Configuration Area Register "RESERVED_3C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AD#) =>
      -- AEB General Configuration Area Register "RESERVED_3CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AE#) =>
      -- AEB General Configuration Area Register "RESERVED_3D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1AF#) =>
      -- AEB General Configuration Area Register "RESERVED_3D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B0#) =>
      -- AEB General Configuration Area Register "RESERVED_3D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B1#) =>
      -- AEB General Configuration Area Register "RESERVED_3DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B2#) =>
      -- AEB General Configuration Area Register "RESERVED_3E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B3#) =>
      -- AEB General Configuration Area Register "RESERVED_3E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B4#) =>
      -- AEB General Configuration Area Register "RESERVED_3E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B5#) =>
      -- AEB General Configuration Area Register "RESERVED_3EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B6#) =>
      -- AEB General Configuration Area Register "RESERVED_3F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B7#) =>
      -- AEB General Configuration Area Register "RESERVED_3F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B8#) =>
      -- AEB General Configuration Area Register "RESERVED_3F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1B9#) =>
      -- AEB General Configuration Area Register "RESERVED_3FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_3fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BA#) =>
      -- AEB General Configuration Area Register "RESERVED_400" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_400.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BB#) =>
      -- AEB General Configuration Area Register "RESERVED_404" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_404.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BC#) =>
      -- AEB General Configuration Area Register "RESERVED_408" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_408.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BD#) =>
      -- AEB General Configuration Area Register "RESERVED_40C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_40c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BE#) =>
      -- AEB General Configuration Area Register "RESERVED_410" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_410.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1BF#) =>
      -- AEB General Configuration Area Register "RESERVED_414" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_414.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C0#) =>
      -- AEB General Configuration Area Register "RESERVED_418" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_418.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C1#) =>
      -- AEB General Configuration Area Register "RESERVED_41C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_41c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C2#) =>
      -- AEB General Configuration Area Register "RESERVED_420" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_420.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C3#) =>
      -- AEB General Configuration Area Register "RESERVED_424" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_424.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C4#) =>
      -- AEB General Configuration Area Register "RESERVED_428" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_428.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C5#) =>
      -- AEB General Configuration Area Register "RESERVED_42C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_42c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C6#) =>
      -- AEB General Configuration Area Register "RESERVED_430" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_430.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C7#) =>
      -- AEB General Configuration Area Register "RESERVED_434" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_434.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C8#) =>
      -- AEB General Configuration Area Register "RESERVED_438" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_438.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1C9#) =>
      -- AEB General Configuration Area Register "RESERVED_43C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_43c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CA#) =>
      -- AEB General Configuration Area Register "RESERVED_440" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_440.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CB#) =>
      -- AEB General Configuration Area Register "RESERVED_444" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_444.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CC#) =>
      -- AEB General Configuration Area Register "RESERVED_448" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_448.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CD#) =>
      -- AEB General Configuration Area Register "RESERVED_44C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_44c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CE#) =>
      -- AEB General Configuration Area Register "RESERVED_450" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_450.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1CF#) =>
      -- AEB General Configuration Area Register "RESERVED_454" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_454.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D0#) =>
      -- AEB General Configuration Area Register "RESERVED_458" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_458.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D1#) =>
      -- AEB General Configuration Area Register "RESERVED_45C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_45c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D2#) =>
      -- AEB General Configuration Area Register "RESERVED_460" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_460.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D3#) =>
      -- AEB General Configuration Area Register "RESERVED_464" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_464.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D4#) =>
      -- AEB General Configuration Area Register "RESERVED_468" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_468.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D5#) =>
      -- AEB General Configuration Area Register "RESERVED_46C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_46c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D6#) =>
      -- AEB General Configuration Area Register "RESERVED_470" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_470.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D7#) =>
      -- AEB General Configuration Area Register "RESERVED_474" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_474.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D8#) =>
      -- AEB General Configuration Area Register "RESERVED_478" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_478.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1D9#) =>
      -- AEB General Configuration Area Register "RESERVED_47C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_47c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DA#) =>
      -- AEB General Configuration Area Register "RESERVED_480" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_480.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DB#) =>
      -- AEB General Configuration Area Register "RESERVED_484" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_484.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DC#) =>
      -- AEB General Configuration Area Register "RESERVED_488" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_488.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DD#) =>
      -- AEB General Configuration Area Register "RESERVED_48C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_48c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DE#) =>
      -- AEB General Configuration Area Register "RESERVED_490" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_490.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1DF#) =>
      -- AEB General Configuration Area Register "RESERVED_494" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_494.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E0#) =>
      -- AEB General Configuration Area Register "RESERVED_498" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_498.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E1#) =>
      -- AEB General Configuration Area Register "RESERVED_49C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_49c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E2#) =>
      -- AEB General Configuration Area Register "RESERVED_4A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E3#) =>
      -- AEB General Configuration Area Register "RESERVED_4A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E4#) =>
      -- AEB General Configuration Area Register "RESERVED_4A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E5#) =>
      -- AEB General Configuration Area Register "RESERVED_4AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E6#) =>
      -- AEB General Configuration Area Register "RESERVED_4B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E7#) =>
      -- AEB General Configuration Area Register "RESERVED_4B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E8#) =>
      -- AEB General Configuration Area Register "RESERVED_4B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1E9#) =>
      -- AEB General Configuration Area Register "RESERVED_4BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1EA#) =>
      -- AEB General Configuration Area Register "RESERVED_4C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1EB#) =>
      -- AEB General Configuration Area Register "RESERVED_4C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1EC#) =>
      -- AEB General Configuration Area Register "RESERVED_4C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1ED#) =>
      -- AEB General Configuration Area Register "RESERVED_4CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1EE#) =>
      -- AEB General Configuration Area Register "RESERVED_4D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1EF#) =>
      -- AEB General Configuration Area Register "RESERVED_4D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F0#) =>
      -- AEB General Configuration Area Register "RESERVED_4D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F1#) =>
      -- AEB General Configuration Area Register "RESERVED_4DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F2#) =>
      -- AEB General Configuration Area Register "RESERVED_4E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F3#) =>
      -- AEB General Configuration Area Register "RESERVED_4E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F4#) =>
      -- AEB General Configuration Area Register "RESERVED_4E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F5#) =>
      -- AEB General Configuration Area Register "RESERVED_4EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F6#) =>
      -- AEB General Configuration Area Register "RESERVED_4F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F7#) =>
      -- AEB General Configuration Area Register "RESERVED_4F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F8#) =>
      -- AEB General Configuration Area Register "RESERVED_4F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1F9#) =>
      -- AEB General Configuration Area Register "RESERVED_4FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_4fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FA#) =>
      -- AEB General Configuration Area Register "RESERVED_500" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_500.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FB#) =>
      -- AEB General Configuration Area Register "RESERVED_504" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_504.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FC#) =>
      -- AEB General Configuration Area Register "RESERVED_508" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_508.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FD#) =>
      -- AEB General Configuration Area Register "RESERVED_50C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_50c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FE#) =>
      -- AEB General Configuration Area Register "RESERVED_510" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_510.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#1FF#) =>
      -- AEB General Configuration Area Register "RESERVED_514" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_514.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#200#) =>
      -- AEB General Configuration Area Register "RESERVED_518" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_518.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#201#) =>
      -- AEB General Configuration Area Register "RESERVED_51C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_51c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#202#) =>
      -- AEB General Configuration Area Register "RESERVED_520" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_520.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#203#) =>
      -- AEB General Configuration Area Register "RESERVED_524" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_524.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#204#) =>
      -- AEB General Configuration Area Register "RESERVED_528" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_528.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#205#) =>
      -- AEB General Configuration Area Register "RESERVED_52C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_52c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#206#) =>
      -- AEB General Configuration Area Register "RESERVED_530" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_530.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#207#) =>
      -- AEB General Configuration Area Register "RESERVED_534" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_534.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#208#) =>
      -- AEB General Configuration Area Register "RESERVED_538" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_538.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#209#) =>
      -- AEB General Configuration Area Register "RESERVED_53C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_53c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20A#) =>
      -- AEB General Configuration Area Register "RESERVED_540" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_540.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20B#) =>
      -- AEB General Configuration Area Register "RESERVED_544" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_544.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20C#) =>
      -- AEB General Configuration Area Register "RESERVED_548" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_548.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20D#) =>
      -- AEB General Configuration Area Register "RESERVED_54C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_54c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20E#) =>
      -- AEB General Configuration Area Register "RESERVED_550" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_550.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#20F#) =>
      -- AEB General Configuration Area Register "RESERVED_554" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_554.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#210#) =>
      -- AEB General Configuration Area Register "RESERVED_558" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_558.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#211#) =>
      -- AEB General Configuration Area Register "RESERVED_55C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_55c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#212#) =>
      -- AEB General Configuration Area Register "RESERVED_560" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_560.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#213#) =>
      -- AEB General Configuration Area Register "RESERVED_564" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_564.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#214#) =>
      -- AEB General Configuration Area Register "RESERVED_568" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_568.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#215#) =>
      -- AEB General Configuration Area Register "RESERVED_56C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_56c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#216#) =>
      -- AEB General Configuration Area Register "RESERVED_570" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_570.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#217#) =>
      -- AEB General Configuration Area Register "RESERVED_574" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_574.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#218#) =>
      -- AEB General Configuration Area Register "RESERVED_578" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_578.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#219#) =>
      -- AEB General Configuration Area Register "RESERVED_57C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_57c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21A#) =>
      -- AEB General Configuration Area Register "RESERVED_580" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_580.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21B#) =>
      -- AEB General Configuration Area Register "RESERVED_584" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_584.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21C#) =>
      -- AEB General Configuration Area Register "RESERVED_588" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_588.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21D#) =>
      -- AEB General Configuration Area Register "RESERVED_58C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_58c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21E#) =>
      -- AEB General Configuration Area Register "RESERVED_590" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_590.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#21F#) =>
      -- AEB General Configuration Area Register "RESERVED_594" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_594.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#220#) =>
      -- AEB General Configuration Area Register "RESERVED_598" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_598.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#221#) =>
      -- AEB General Configuration Area Register "RESERVED_59C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_59c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#222#) =>
      -- AEB General Configuration Area Register "RESERVED_5A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#223#) =>
      -- AEB General Configuration Area Register "RESERVED_5A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#224#) =>
      -- AEB General Configuration Area Register "RESERVED_5A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#225#) =>
      -- AEB General Configuration Area Register "RESERVED_5AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#226#) =>
      -- AEB General Configuration Area Register "RESERVED_5B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#227#) =>
      -- AEB General Configuration Area Register "RESERVED_5B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#228#) =>
      -- AEB General Configuration Area Register "RESERVED_5B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#229#) =>
      -- AEB General Configuration Area Register "RESERVED_5BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22A#) =>
      -- AEB General Configuration Area Register "RESERVED_5C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22B#) =>
      -- AEB General Configuration Area Register "RESERVED_5C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22C#) =>
      -- AEB General Configuration Area Register "RESERVED_5C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22D#) =>
      -- AEB General Configuration Area Register "RESERVED_5CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22E#) =>
      -- AEB General Configuration Area Register "RESERVED_5D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#22F#) =>
      -- AEB General Configuration Area Register "RESERVED_5D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#230#) =>
      -- AEB General Configuration Area Register "RESERVED_5D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#231#) =>
      -- AEB General Configuration Area Register "RESERVED_5DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#232#) =>
      -- AEB General Configuration Area Register "RESERVED_5E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#233#) =>
      -- AEB General Configuration Area Register "RESERVED_5E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#234#) =>
      -- AEB General Configuration Area Register "RESERVED_5E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#235#) =>
      -- AEB General Configuration Area Register "RESERVED_5EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#236#) =>
      -- AEB General Configuration Area Register "RESERVED_5F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#237#) =>
      -- AEB General Configuration Area Register "RESERVED_5F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#238#) =>
      -- AEB General Configuration Area Register "RESERVED_5F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#239#) =>
      -- AEB General Configuration Area Register "RESERVED_5FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_5fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23A#) =>
      -- AEB General Configuration Area Register "RESERVED_600" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_600.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23B#) =>
      -- AEB General Configuration Area Register "RESERVED_604" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_604.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23C#) =>
      -- AEB General Configuration Area Register "RESERVED_608" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_608.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23D#) =>
      -- AEB General Configuration Area Register "RESERVED_60C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_60c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23E#) =>
      -- AEB General Configuration Area Register "RESERVED_610" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_610.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#23F#) =>
      -- AEB General Configuration Area Register "RESERVED_614" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_614.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#240#) =>
      -- AEB General Configuration Area Register "RESERVED_618" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_618.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#241#) =>
      -- AEB General Configuration Area Register "RESERVED_61C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_61c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#242#) =>
      -- AEB General Configuration Area Register "RESERVED_620" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_620.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#243#) =>
      -- AEB General Configuration Area Register "RESERVED_624" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_624.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#244#) =>
      -- AEB General Configuration Area Register "RESERVED_628" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_628.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#245#) =>
      -- AEB General Configuration Area Register "RESERVED_62C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_62c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#246#) =>
      -- AEB General Configuration Area Register "RESERVED_630" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_630.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#247#) =>
      -- AEB General Configuration Area Register "RESERVED_634" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_634.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#248#) =>
      -- AEB General Configuration Area Register "RESERVED_638" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_638.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#249#) =>
      -- AEB General Configuration Area Register "RESERVED_63C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_63c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24A#) =>
      -- AEB General Configuration Area Register "RESERVED_640" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_640.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24B#) =>
      -- AEB General Configuration Area Register "RESERVED_644" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_644.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24C#) =>
      -- AEB General Configuration Area Register "RESERVED_648" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_648.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24D#) =>
      -- AEB General Configuration Area Register "RESERVED_64C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_64c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24E#) =>
      -- AEB General Configuration Area Register "RESERVED_650" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_650.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#24F#) =>
      -- AEB General Configuration Area Register "RESERVED_654" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_654.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#250#) =>
      -- AEB General Configuration Area Register "RESERVED_658" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_658.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#251#) =>
      -- AEB General Configuration Area Register "RESERVED_65C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_65c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#252#) =>
      -- AEB General Configuration Area Register "RESERVED_660" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_660.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#253#) =>
      -- AEB General Configuration Area Register "RESERVED_664" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_664.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#254#) =>
      -- AEB General Configuration Area Register "RESERVED_668" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_668.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#255#) =>
      -- AEB General Configuration Area Register "RESERVED_66C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_66c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#256#) =>
      -- AEB General Configuration Area Register "RESERVED_670" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_670.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#257#) =>
      -- AEB General Configuration Area Register "RESERVED_674" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_674.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#258#) =>
      -- AEB General Configuration Area Register "RESERVED_678" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_678.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#259#) =>
      -- AEB General Configuration Area Register "RESERVED_67C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_67c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25A#) =>
      -- AEB General Configuration Area Register "RESERVED_680" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_680.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25B#) =>
      -- AEB General Configuration Area Register "RESERVED_684" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_684.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25C#) =>
      -- AEB General Configuration Area Register "RESERVED_688" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_688.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25D#) =>
      -- AEB General Configuration Area Register "RESERVED_68C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_68c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25E#) =>
      -- AEB General Configuration Area Register "RESERVED_690" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_690.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#25F#) =>
      -- AEB General Configuration Area Register "RESERVED_694" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_694.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#260#) =>
      -- AEB General Configuration Area Register "RESERVED_698" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_698.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#261#) =>
      -- AEB General Configuration Area Register "RESERVED_69C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_69c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#262#) =>
      -- AEB General Configuration Area Register "RESERVED_6A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#263#) =>
      -- AEB General Configuration Area Register "RESERVED_6A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#264#) =>
      -- AEB General Configuration Area Register "RESERVED_6A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#265#) =>
      -- AEB General Configuration Area Register "RESERVED_6AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#266#) =>
      -- AEB General Configuration Area Register "RESERVED_6B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#267#) =>
      -- AEB General Configuration Area Register "RESERVED_6B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#268#) =>
      -- AEB General Configuration Area Register "RESERVED_6B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#269#) =>
      -- AEB General Configuration Area Register "RESERVED_6BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26A#) =>
      -- AEB General Configuration Area Register "RESERVED_6C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26B#) =>
      -- AEB General Configuration Area Register "RESERVED_6C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26C#) =>
      -- AEB General Configuration Area Register "RESERVED_6C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26D#) =>
      -- AEB General Configuration Area Register "RESERVED_6CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26E#) =>
      -- AEB General Configuration Area Register "RESERVED_6D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#26F#) =>
      -- AEB General Configuration Area Register "RESERVED_6D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#270#) =>
      -- AEB General Configuration Area Register "RESERVED_6D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#271#) =>
      -- AEB General Configuration Area Register "RESERVED_6DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#272#) =>
      -- AEB General Configuration Area Register "RESERVED_6E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#273#) =>
      -- AEB General Configuration Area Register "RESERVED_6E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#274#) =>
      -- AEB General Configuration Area Register "RESERVED_6E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#275#) =>
      -- AEB General Configuration Area Register "RESERVED_6EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#276#) =>
      -- AEB General Configuration Area Register "RESERVED_6F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#277#) =>
      -- AEB General Configuration Area Register "RESERVED_6F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#278#) =>
      -- AEB General Configuration Area Register "RESERVED_6F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#279#) =>
      -- AEB General Configuration Area Register "RESERVED_6FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_6fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27A#) =>
      -- AEB General Configuration Area Register "RESERVED_700" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_700.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27B#) =>
      -- AEB General Configuration Area Register "RESERVED_704" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_704.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27C#) =>
      -- AEB General Configuration Area Register "RESERVED_708" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_708.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27D#) =>
      -- AEB General Configuration Area Register "RESERVED_70C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_70c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27E#) =>
      -- AEB General Configuration Area Register "RESERVED_710" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_710.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#27F#) =>
      -- AEB General Configuration Area Register "RESERVED_714" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_714.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#280#) =>
      -- AEB General Configuration Area Register "RESERVED_718" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_718.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#281#) =>
      -- AEB General Configuration Area Register "RESERVED_71C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_71c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#282#) =>
      -- AEB General Configuration Area Register "RESERVED_720" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_720.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#283#) =>
      -- AEB General Configuration Area Register "RESERVED_724" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_724.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#284#) =>
      -- AEB General Configuration Area Register "RESERVED_728" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_728.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#285#) =>
      -- AEB General Configuration Area Register "RESERVED_72C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_72c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#286#) =>
      -- AEB General Configuration Area Register "RESERVED_730" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_730.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#287#) =>
      -- AEB General Configuration Area Register "RESERVED_734" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_734.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#288#) =>
      -- AEB General Configuration Area Register "RESERVED_738" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_738.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#289#) =>
      -- AEB General Configuration Area Register "RESERVED_73C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_73c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28A#) =>
      -- AEB General Configuration Area Register "RESERVED_740" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_740.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28B#) =>
      -- AEB General Configuration Area Register "RESERVED_744" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_744.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28C#) =>
      -- AEB General Configuration Area Register "RESERVED_748" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_748.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28D#) =>
      -- AEB General Configuration Area Register "RESERVED_74C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_74c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28E#) =>
      -- AEB General Configuration Area Register "RESERVED_750" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_750.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#28F#) =>
      -- AEB General Configuration Area Register "RESERVED_754" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_754.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#290#) =>
      -- AEB General Configuration Area Register "RESERVED_758" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_758.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#291#) =>
      -- AEB General Configuration Area Register "RESERVED_75C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_75c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#292#) =>
      -- AEB General Configuration Area Register "RESERVED_760" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_760.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#293#) =>
      -- AEB General Configuration Area Register "RESERVED_764" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_764.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#294#) =>
      -- AEB General Configuration Area Register "RESERVED_768" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_768.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#295#) =>
      -- AEB General Configuration Area Register "RESERVED_76C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_76c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#296#) =>
      -- AEB General Configuration Area Register "RESERVED_770" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_770.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#297#) =>
      -- AEB General Configuration Area Register "RESERVED_774" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_774.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#298#) =>
      -- AEB General Configuration Area Register "RESERVED_778" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_778.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#299#) =>
      -- AEB General Configuration Area Register "RESERVED_77C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_77c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29A#) =>
      -- AEB General Configuration Area Register "RESERVED_780" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_780.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29B#) =>
      -- AEB General Configuration Area Register "RESERVED_784" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_784.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29C#) =>
      -- AEB General Configuration Area Register "RESERVED_788" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_788.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29D#) =>
      -- AEB General Configuration Area Register "RESERVED_78C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_78c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29E#) =>
      -- AEB General Configuration Area Register "RESERVED_790" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_790.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#29F#) =>
      -- AEB General Configuration Area Register "RESERVED_794" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_794.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A0#) =>
      -- AEB General Configuration Area Register "RESERVED_798" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_798.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A1#) =>
      -- AEB General Configuration Area Register "RESERVED_79C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_79c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A2#) =>
      -- AEB General Configuration Area Register "RESERVED_7A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A3#) =>
      -- AEB General Configuration Area Register "RESERVED_7A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A4#) =>
      -- AEB General Configuration Area Register "RESERVED_7A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A5#) =>
      -- AEB General Configuration Area Register "RESERVED_7AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A6#) =>
      -- AEB General Configuration Area Register "RESERVED_7B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A7#) =>
      -- AEB General Configuration Area Register "RESERVED_7B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A8#) =>
      -- AEB General Configuration Area Register "RESERVED_7B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2A9#) =>
      -- AEB General Configuration Area Register "RESERVED_7BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AA#) =>
      -- AEB General Configuration Area Register "RESERVED_7C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AB#) =>
      -- AEB General Configuration Area Register "RESERVED_7C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AC#) =>
      -- AEB General Configuration Area Register "RESERVED_7C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AD#) =>
      -- AEB General Configuration Area Register "RESERVED_7CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AE#) =>
      -- AEB General Configuration Area Register "RESERVED_7D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2AF#) =>
      -- AEB General Configuration Area Register "RESERVED_7D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B0#) =>
      -- AEB General Configuration Area Register "RESERVED_7D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B1#) =>
      -- AEB General Configuration Area Register "RESERVED_7DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B2#) =>
      -- AEB General Configuration Area Register "RESERVED_7E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B3#) =>
      -- AEB General Configuration Area Register "RESERVED_7E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B4#) =>
      -- AEB General Configuration Area Register "RESERVED_7E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B5#) =>
      -- AEB General Configuration Area Register "RESERVED_7EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B6#) =>
      -- AEB General Configuration Area Register "RESERVED_7F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B7#) =>
      -- AEB General Configuration Area Register "RESERVED_7F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B8#) =>
      -- AEB General Configuration Area Register "RESERVED_7F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2B9#) =>
      -- AEB General Configuration Area Register "RESERVED_7FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_7fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BA#) =>
      -- AEB General Configuration Area Register "RESERVED_800" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_800.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BB#) =>
      -- AEB General Configuration Area Register "RESERVED_804" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_804.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BC#) =>
      -- AEB General Configuration Area Register "RESERVED_808" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_808.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BD#) =>
      -- AEB General Configuration Area Register "RESERVED_80C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_80c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BE#) =>
      -- AEB General Configuration Area Register "RESERVED_810" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_810.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2BF#) =>
      -- AEB General Configuration Area Register "RESERVED_814" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_814.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C0#) =>
      -- AEB General Configuration Area Register "RESERVED_818" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_818.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C1#) =>
      -- AEB General Configuration Area Register "RESERVED_81C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_81c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C2#) =>
      -- AEB General Configuration Area Register "RESERVED_820" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_820.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C3#) =>
      -- AEB General Configuration Area Register "RESERVED_824" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_824.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C4#) =>
      -- AEB General Configuration Area Register "RESERVED_828" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_828.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C5#) =>
      -- AEB General Configuration Area Register "RESERVED_82C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_82c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C6#) =>
      -- AEB General Configuration Area Register "RESERVED_830" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_830.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C7#) =>
      -- AEB General Configuration Area Register "RESERVED_834" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_834.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C8#) =>
      -- AEB General Configuration Area Register "RESERVED_838" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_838.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2C9#) =>
      -- AEB General Configuration Area Register "RESERVED_83C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_83c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CA#) =>
      -- AEB General Configuration Area Register "RESERVED_840" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_840.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CB#) =>
      -- AEB General Configuration Area Register "RESERVED_844" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_844.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CC#) =>
      -- AEB General Configuration Area Register "RESERVED_848" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_848.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CD#) =>
      -- AEB General Configuration Area Register "RESERVED_84C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_84c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CE#) =>
      -- AEB General Configuration Area Register "RESERVED_850" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_850.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2CF#) =>
      -- AEB General Configuration Area Register "RESERVED_854" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_854.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D0#) =>
      -- AEB General Configuration Area Register "RESERVED_858" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_858.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D1#) =>
      -- AEB General Configuration Area Register "RESERVED_85C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_85c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D2#) =>
      -- AEB General Configuration Area Register "RESERVED_860" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_860.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D3#) =>
      -- AEB General Configuration Area Register "RESERVED_864" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_864.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D4#) =>
      -- AEB General Configuration Area Register "RESERVED_868" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_868.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D5#) =>
      -- AEB General Configuration Area Register "RESERVED_86C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_86c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D6#) =>
      -- AEB General Configuration Area Register "RESERVED_870" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_870.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D7#) =>
      -- AEB General Configuration Area Register "RESERVED_874" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_874.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D8#) =>
      -- AEB General Configuration Area Register "RESERVED_878" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_878.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2D9#) =>
      -- AEB General Configuration Area Register "RESERVED_87C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_87c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DA#) =>
      -- AEB General Configuration Area Register "RESERVED_880" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_880.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DB#) =>
      -- AEB General Configuration Area Register "RESERVED_884" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_884.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DC#) =>
      -- AEB General Configuration Area Register "RESERVED_888" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_888.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DD#) =>
      -- AEB General Configuration Area Register "RESERVED_88C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_88c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DE#) =>
      -- AEB General Configuration Area Register "RESERVED_890" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_890.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2DF#) =>
      -- AEB General Configuration Area Register "RESERVED_894" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_894.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E0#) =>
      -- AEB General Configuration Area Register "RESERVED_898" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_898.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E1#) =>
      -- AEB General Configuration Area Register "RESERVED_89C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_89c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E2#) =>
      -- AEB General Configuration Area Register "RESERVED_8A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E3#) =>
      -- AEB General Configuration Area Register "RESERVED_8A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E4#) =>
      -- AEB General Configuration Area Register "RESERVED_8A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E5#) =>
      -- AEB General Configuration Area Register "RESERVED_8AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E6#) =>
      -- AEB General Configuration Area Register "RESERVED_8B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E7#) =>
      -- AEB General Configuration Area Register "RESERVED_8B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E8#) =>
      -- AEB General Configuration Area Register "RESERVED_8B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2E9#) =>
      -- AEB General Configuration Area Register "RESERVED_8BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2EA#) =>
      -- AEB General Configuration Area Register "RESERVED_8C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2EB#) =>
      -- AEB General Configuration Area Register "RESERVED_8C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2EC#) =>
      -- AEB General Configuration Area Register "RESERVED_8C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2ED#) =>
      -- AEB General Configuration Area Register "RESERVED_8CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2EE#) =>
      -- AEB General Configuration Area Register "RESERVED_8D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2EF#) =>
      -- AEB General Configuration Area Register "RESERVED_8D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F0#) =>
      -- AEB General Configuration Area Register "RESERVED_8D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F1#) =>
      -- AEB General Configuration Area Register "RESERVED_8DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F2#) =>
      -- AEB General Configuration Area Register "RESERVED_8E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F3#) =>
      -- AEB General Configuration Area Register "RESERVED_8E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F4#) =>
      -- AEB General Configuration Area Register "RESERVED_8E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F5#) =>
      -- AEB General Configuration Area Register "RESERVED_8EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F6#) =>
      -- AEB General Configuration Area Register "RESERVED_8F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F7#) =>
      -- AEB General Configuration Area Register "RESERVED_8F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F8#) =>
      -- AEB General Configuration Area Register "RESERVED_8F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2F9#) =>
      -- AEB General Configuration Area Register "RESERVED_8FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_8fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FA#) =>
      -- AEB General Configuration Area Register "RESERVED_900" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_900.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FB#) =>
      -- AEB General Configuration Area Register "RESERVED_904" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_904.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FC#) =>
      -- AEB General Configuration Area Register "RESERVED_908" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_908.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FD#) =>
      -- AEB General Configuration Area Register "RESERVED_90C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_90c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FE#) =>
      -- AEB General Configuration Area Register "RESERVED_910" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_910.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#2FF#) =>
      -- AEB General Configuration Area Register "RESERVED_914" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_914.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#300#) =>
      -- AEB General Configuration Area Register "RESERVED_918" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_918.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#301#) =>
      -- AEB General Configuration Area Register "RESERVED_91C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_91c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#302#) =>
      -- AEB General Configuration Area Register "RESERVED_920" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_920.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#303#) =>
      -- AEB General Configuration Area Register "RESERVED_924" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_924.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#304#) =>
      -- AEB General Configuration Area Register "RESERVED_928" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_928.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#305#) =>
      -- AEB General Configuration Area Register "RESERVED_92C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_92c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#306#) =>
      -- AEB General Configuration Area Register "RESERVED_930" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_930.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#307#) =>
      -- AEB General Configuration Area Register "RESERVED_934" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_934.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#308#) =>
      -- AEB General Configuration Area Register "RESERVED_938" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_938.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#309#) =>
      -- AEB General Configuration Area Register "RESERVED_93C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_93c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30A#) =>
      -- AEB General Configuration Area Register "RESERVED_940" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_940.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30B#) =>
      -- AEB General Configuration Area Register "RESERVED_944" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_944.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30C#) =>
      -- AEB General Configuration Area Register "RESERVED_948" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_948.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30D#) =>
      -- AEB General Configuration Area Register "RESERVED_94C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_94c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30E#) =>
      -- AEB General Configuration Area Register "RESERVED_950" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_950.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#30F#) =>
      -- AEB General Configuration Area Register "RESERVED_954" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_954.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#310#) =>
      -- AEB General Configuration Area Register "RESERVED_958" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_958.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#311#) =>
      -- AEB General Configuration Area Register "RESERVED_95C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_95c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#312#) =>
      -- AEB General Configuration Area Register "RESERVED_960" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_960.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#313#) =>
      -- AEB General Configuration Area Register "RESERVED_964" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_964.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#314#) =>
      -- AEB General Configuration Area Register "RESERVED_968" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_968.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#315#) =>
      -- AEB General Configuration Area Register "RESERVED_96C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_96c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#316#) =>
      -- AEB General Configuration Area Register "RESERVED_970" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_970.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#317#) =>
      -- AEB General Configuration Area Register "RESERVED_974" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_974.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#318#) =>
      -- AEB General Configuration Area Register "RESERVED_978" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_978.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#319#) =>
      -- AEB General Configuration Area Register "RESERVED_97C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_97c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31A#) =>
      -- AEB General Configuration Area Register "RESERVED_980" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_980.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31B#) =>
      -- AEB General Configuration Area Register "RESERVED_984" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_984.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31C#) =>
      -- AEB General Configuration Area Register "RESERVED_988" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_988.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31D#) =>
      -- AEB General Configuration Area Register "RESERVED_98C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_98c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31E#) =>
      -- AEB General Configuration Area Register "RESERVED_990" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_990.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#31F#) =>
      -- AEB General Configuration Area Register "RESERVED_994" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_994.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#320#) =>
      -- AEB General Configuration Area Register "RESERVED_998" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_998.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#321#) =>
      -- AEB General Configuration Area Register "RESERVED_99C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_99c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#322#) =>
      -- AEB General Configuration Area Register "RESERVED_9A0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#323#) =>
      -- AEB General Configuration Area Register "RESERVED_9A4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#324#) =>
      -- AEB General Configuration Area Register "RESERVED_9A8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9a8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#325#) =>
      -- AEB General Configuration Area Register "RESERVED_9AC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#326#) =>
      -- AEB General Configuration Area Register "RESERVED_9B0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#327#) =>
      -- AEB General Configuration Area Register "RESERVED_9B4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#328#) =>
      -- AEB General Configuration Area Register "RESERVED_9B8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9b8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#329#) =>
      -- AEB General Configuration Area Register "RESERVED_9BC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9bc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32A#) =>
      -- AEB General Configuration Area Register "RESERVED_9C0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32B#) =>
      -- AEB General Configuration Area Register "RESERVED_9C4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32C#) =>
      -- AEB General Configuration Area Register "RESERVED_9C8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9c8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32D#) =>
      -- AEB General Configuration Area Register "RESERVED_9CC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9cc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32E#) =>
      -- AEB General Configuration Area Register "RESERVED_9D0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#32F#) =>
      -- AEB General Configuration Area Register "RESERVED_9D4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#330#) =>
      -- AEB General Configuration Area Register "RESERVED_9D8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9d8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#331#) =>
      -- AEB General Configuration Area Register "RESERVED_9DC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9dc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#332#) =>
      -- AEB General Configuration Area Register "RESERVED_9E0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#333#) =>
      -- AEB General Configuration Area Register "RESERVED_9E4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#334#) =>
      -- AEB General Configuration Area Register "RESERVED_9E8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9e8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#335#) =>
      -- AEB General Configuration Area Register "RESERVED_9EC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9ec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#336#) =>
      -- AEB General Configuration Area Register "RESERVED_9F0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#337#) =>
      -- AEB General Configuration Area Register "RESERVED_9F4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#338#) =>
      -- AEB General Configuration Area Register "RESERVED_9F8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9f8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#339#) =>
      -- AEB General Configuration Area Register "RESERVED_9FC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_9fc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33A#) =>
      -- AEB General Configuration Area Register "RESERVED_A00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33B#) =>
      -- AEB General Configuration Area Register "RESERVED_A04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33C#) =>
      -- AEB General Configuration Area Register "RESERVED_A08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33D#) =>
      -- AEB General Configuration Area Register "RESERVED_A0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33E#) =>
      -- AEB General Configuration Area Register "RESERVED_A10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#33F#) =>
      -- AEB General Configuration Area Register "RESERVED_A14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#340#) =>
      -- AEB General Configuration Area Register "RESERVED_A18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#341#) =>
      -- AEB General Configuration Area Register "RESERVED_A1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#342#) =>
      -- AEB General Configuration Area Register "RESERVED_A20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#343#) =>
      -- AEB General Configuration Area Register "RESERVED_A24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#344#) =>
      -- AEB General Configuration Area Register "RESERVED_A28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#345#) =>
      -- AEB General Configuration Area Register "RESERVED_A2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#346#) =>
      -- AEB General Configuration Area Register "RESERVED_A30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#347#) =>
      -- AEB General Configuration Area Register "RESERVED_A34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#348#) =>
      -- AEB General Configuration Area Register "RESERVED_A38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#349#) =>
      -- AEB General Configuration Area Register "RESERVED_A3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34A#) =>
      -- AEB General Configuration Area Register "RESERVED_A40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34B#) =>
      -- AEB General Configuration Area Register "RESERVED_A44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34C#) =>
      -- AEB General Configuration Area Register "RESERVED_A48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34D#) =>
      -- AEB General Configuration Area Register "RESERVED_A4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34E#) =>
      -- AEB General Configuration Area Register "RESERVED_A50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#34F#) =>
      -- AEB General Configuration Area Register "RESERVED_A54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#350#) =>
      -- AEB General Configuration Area Register "RESERVED_A58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#351#) =>
      -- AEB General Configuration Area Register "RESERVED_A5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#352#) =>
      -- AEB General Configuration Area Register "RESERVED_A60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#353#) =>
      -- AEB General Configuration Area Register "RESERVED_A64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#354#) =>
      -- AEB General Configuration Area Register "RESERVED_A68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#355#) =>
      -- AEB General Configuration Area Register "RESERVED_A6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#356#) =>
      -- AEB General Configuration Area Register "RESERVED_A70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#357#) =>
      -- AEB General Configuration Area Register "RESERVED_A74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#358#) =>
      -- AEB General Configuration Area Register "RESERVED_A78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#359#) =>
      -- AEB General Configuration Area Register "RESERVED_A7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35A#) =>
      -- AEB General Configuration Area Register "RESERVED_A80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35B#) =>
      -- AEB General Configuration Area Register "RESERVED_A84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35C#) =>
      -- AEB General Configuration Area Register "RESERVED_A88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35D#) =>
      -- AEB General Configuration Area Register "RESERVED_A8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35E#) =>
      -- AEB General Configuration Area Register "RESERVED_A90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#35F#) =>
      -- AEB General Configuration Area Register "RESERVED_A94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#360#) =>
      -- AEB General Configuration Area Register "RESERVED_A98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#361#) =>
      -- AEB General Configuration Area Register "RESERVED_A9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_a9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#362#) =>
      -- AEB General Configuration Area Register "RESERVED_AA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#363#) =>
      -- AEB General Configuration Area Register "RESERVED_AA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#364#) =>
      -- AEB General Configuration Area Register "RESERVED_AA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aa8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#365#) =>
      -- AEB General Configuration Area Register "RESERVED_AAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#366#) =>
      -- AEB General Configuration Area Register "RESERVED_AB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#367#) =>
      -- AEB General Configuration Area Register "RESERVED_AB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#368#) =>
      -- AEB General Configuration Area Register "RESERVED_AB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ab8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#369#) =>
      -- AEB General Configuration Area Register "RESERVED_ABC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_abc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36A#) =>
      -- AEB General Configuration Area Register "RESERVED_AC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36B#) =>
      -- AEB General Configuration Area Register "RESERVED_AC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36C#) =>
      -- AEB General Configuration Area Register "RESERVED_AC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ac8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36D#) =>
      -- AEB General Configuration Area Register "RESERVED_ACC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_acc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36E#) =>
      -- AEB General Configuration Area Register "RESERVED_AD0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#36F#) =>
      -- AEB General Configuration Area Register "RESERVED_AD4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#370#) =>
      -- AEB General Configuration Area Register "RESERVED_AD8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ad8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#371#) =>
      -- AEB General Configuration Area Register "RESERVED_ADC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_adc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#372#) =>
      -- AEB General Configuration Area Register "RESERVED_AE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#373#) =>
      -- AEB General Configuration Area Register "RESERVED_AE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#374#) =>
      -- AEB General Configuration Area Register "RESERVED_AE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ae8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#375#) =>
      -- AEB General Configuration Area Register "RESERVED_AEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_aec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#376#) =>
      -- AEB General Configuration Area Register "RESERVED_AF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#377#) =>
      -- AEB General Configuration Area Register "RESERVED_AF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#378#) =>
      -- AEB General Configuration Area Register "RESERVED_AF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_af8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#379#) =>
      -- AEB General Configuration Area Register "RESERVED_AFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_afc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37A#) =>
      -- AEB General Configuration Area Register "RESERVED_B00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37B#) =>
      -- AEB General Configuration Area Register "RESERVED_B04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37C#) =>
      -- AEB General Configuration Area Register "RESERVED_B08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37D#) =>
      -- AEB General Configuration Area Register "RESERVED_B0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37E#) =>
      -- AEB General Configuration Area Register "RESERVED_B10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#37F#) =>
      -- AEB General Configuration Area Register "RESERVED_B14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#380#) =>
      -- AEB General Configuration Area Register "RESERVED_B18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#381#) =>
      -- AEB General Configuration Area Register "RESERVED_B1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#382#) =>
      -- AEB General Configuration Area Register "RESERVED_B20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#383#) =>
      -- AEB General Configuration Area Register "RESERVED_B24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#384#) =>
      -- AEB General Configuration Area Register "RESERVED_B28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#385#) =>
      -- AEB General Configuration Area Register "RESERVED_B2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#386#) =>
      -- AEB General Configuration Area Register "RESERVED_B30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#387#) =>
      -- AEB General Configuration Area Register "RESERVED_B34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#388#) =>
      -- AEB General Configuration Area Register "RESERVED_B38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#389#) =>
      -- AEB General Configuration Area Register "RESERVED_B3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38A#) =>
      -- AEB General Configuration Area Register "RESERVED_B40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38B#) =>
      -- AEB General Configuration Area Register "RESERVED_B44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38C#) =>
      -- AEB General Configuration Area Register "RESERVED_B48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38D#) =>
      -- AEB General Configuration Area Register "RESERVED_B4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38E#) =>
      -- AEB General Configuration Area Register "RESERVED_B50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#38F#) =>
      -- AEB General Configuration Area Register "RESERVED_B54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#390#) =>
      -- AEB General Configuration Area Register "RESERVED_B58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#391#) =>
      -- AEB General Configuration Area Register "RESERVED_B5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#392#) =>
      -- AEB General Configuration Area Register "RESERVED_B60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#393#) =>
      -- AEB General Configuration Area Register "RESERVED_B64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#394#) =>
      -- AEB General Configuration Area Register "RESERVED_B68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#395#) =>
      -- AEB General Configuration Area Register "RESERVED_B6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#396#) =>
      -- AEB General Configuration Area Register "RESERVED_B70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#397#) =>
      -- AEB General Configuration Area Register "RESERVED_B74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#398#) =>
      -- AEB General Configuration Area Register "RESERVED_B78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#399#) =>
      -- AEB General Configuration Area Register "RESERVED_B7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39A#) =>
      -- AEB General Configuration Area Register "RESERVED_B80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39B#) =>
      -- AEB General Configuration Area Register "RESERVED_B84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39C#) =>
      -- AEB General Configuration Area Register "RESERVED_B88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39D#) =>
      -- AEB General Configuration Area Register "RESERVED_B8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39E#) =>
      -- AEB General Configuration Area Register "RESERVED_B90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#39F#) =>
      -- AEB General Configuration Area Register "RESERVED_B94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A0#) =>
      -- AEB General Configuration Area Register "RESERVED_B98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A1#) =>
      -- AEB General Configuration Area Register "RESERVED_B9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_b9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A2#) =>
      -- AEB General Configuration Area Register "RESERVED_BA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A3#) =>
      -- AEB General Configuration Area Register "RESERVED_BA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A4#) =>
      -- AEB General Configuration Area Register "RESERVED_BA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ba8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A5#) =>
      -- AEB General Configuration Area Register "RESERVED_BAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A6#) =>
      -- AEB General Configuration Area Register "RESERVED_BB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A7#) =>
      -- AEB General Configuration Area Register "RESERVED_BB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A8#) =>
      -- AEB General Configuration Area Register "RESERVED_BB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bb8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3A9#) =>
      -- AEB General Configuration Area Register "RESERVED_BBC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bbc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AA#) =>
      -- AEB General Configuration Area Register "RESERVED_BC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AB#) =>
      -- AEB General Configuration Area Register "RESERVED_BC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AC#) =>
      -- AEB General Configuration Area Register "RESERVED_BC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bc8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AD#) =>
      -- AEB General Configuration Area Register "RESERVED_BCC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bcc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AE#) =>
      -- AEB General Configuration Area Register "RESERVED_BD0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3AF#) =>
      -- AEB General Configuration Area Register "RESERVED_BD4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B0#) =>
      -- AEB General Configuration Area Register "RESERVED_BD8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bd8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B1#) =>
      -- AEB General Configuration Area Register "RESERVED_BDC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bdc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B2#) =>
      -- AEB General Configuration Area Register "RESERVED_BE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B3#) =>
      -- AEB General Configuration Area Register "RESERVED_BE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B4#) =>
      -- AEB General Configuration Area Register "RESERVED_BE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_be8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B5#) =>
      -- AEB General Configuration Area Register "RESERVED_BEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B6#) =>
      -- AEB General Configuration Area Register "RESERVED_BF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B7#) =>
      -- AEB General Configuration Area Register "RESERVED_BF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B8#) =>
      -- AEB General Configuration Area Register "RESERVED_BF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bf8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3B9#) =>
      -- AEB General Configuration Area Register "RESERVED_BFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_bfc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BA#) =>
      -- AEB General Configuration Area Register "RESERVED_C00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BB#) =>
      -- AEB General Configuration Area Register "RESERVED_C04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BC#) =>
      -- AEB General Configuration Area Register "RESERVED_C08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BD#) =>
      -- AEB General Configuration Area Register "RESERVED_C0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BE#) =>
      -- AEB General Configuration Area Register "RESERVED_C10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3BF#) =>
      -- AEB General Configuration Area Register "RESERVED_C14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C0#) =>
      -- AEB General Configuration Area Register "RESERVED_C18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C1#) =>
      -- AEB General Configuration Area Register "RESERVED_C1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C2#) =>
      -- AEB General Configuration Area Register "RESERVED_C20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C3#) =>
      -- AEB General Configuration Area Register "RESERVED_C24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C4#) =>
      -- AEB General Configuration Area Register "RESERVED_C28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C5#) =>
      -- AEB General Configuration Area Register "RESERVED_C2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C6#) =>
      -- AEB General Configuration Area Register "RESERVED_C30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C7#) =>
      -- AEB General Configuration Area Register "RESERVED_C34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C8#) =>
      -- AEB General Configuration Area Register "RESERVED_C38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3C9#) =>
      -- AEB General Configuration Area Register "RESERVED_C3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CA#) =>
      -- AEB General Configuration Area Register "RESERVED_C40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CB#) =>
      -- AEB General Configuration Area Register "RESERVED_C44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CC#) =>
      -- AEB General Configuration Area Register "RESERVED_C48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CD#) =>
      -- AEB General Configuration Area Register "RESERVED_C4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CE#) =>
      -- AEB General Configuration Area Register "RESERVED_C50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3CF#) =>
      -- AEB General Configuration Area Register "RESERVED_C54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D0#) =>
      -- AEB General Configuration Area Register "RESERVED_C58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D1#) =>
      -- AEB General Configuration Area Register "RESERVED_C5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D2#) =>
      -- AEB General Configuration Area Register "RESERVED_C60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D3#) =>
      -- AEB General Configuration Area Register "RESERVED_C64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D4#) =>
      -- AEB General Configuration Area Register "RESERVED_C68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D5#) =>
      -- AEB General Configuration Area Register "RESERVED_C6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D6#) =>
      -- AEB General Configuration Area Register "RESERVED_C70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D7#) =>
      -- AEB General Configuration Area Register "RESERVED_C74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D8#) =>
      -- AEB General Configuration Area Register "RESERVED_C78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3D9#) =>
      -- AEB General Configuration Area Register "RESERVED_C7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DA#) =>
      -- AEB General Configuration Area Register "RESERVED_C80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DB#) =>
      -- AEB General Configuration Area Register "RESERVED_C84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DC#) =>
      -- AEB General Configuration Area Register "RESERVED_C88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DD#) =>
      -- AEB General Configuration Area Register "RESERVED_C8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DE#) =>
      -- AEB General Configuration Area Register "RESERVED_C90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3DF#) =>
      -- AEB General Configuration Area Register "RESERVED_C94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E0#) =>
      -- AEB General Configuration Area Register "RESERVED_C98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E1#) =>
      -- AEB General Configuration Area Register "RESERVED_C9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_c9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E2#) =>
      -- AEB General Configuration Area Register "RESERVED_CA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E3#) =>
      -- AEB General Configuration Area Register "RESERVED_CA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E4#) =>
      -- AEB General Configuration Area Register "RESERVED_CA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ca8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E5#) =>
      -- AEB General Configuration Area Register "RESERVED_CAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E6#) =>
      -- AEB General Configuration Area Register "RESERVED_CB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E7#) =>
      -- AEB General Configuration Area Register "RESERVED_CB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E8#) =>
      -- AEB General Configuration Area Register "RESERVED_CB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cb8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3E9#) =>
      -- AEB General Configuration Area Register "RESERVED_CBC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cbc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3EA#) =>
      -- AEB General Configuration Area Register "RESERVED_CC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3EB#) =>
      -- AEB General Configuration Area Register "RESERVED_CC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3EC#) =>
      -- AEB General Configuration Area Register "RESERVED_CC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cc8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3ED#) =>
      -- AEB General Configuration Area Register "RESERVED_CCC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ccc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3EE#) =>
      -- AEB General Configuration Area Register "RESERVED_CD0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3EF#) =>
      -- AEB General Configuration Area Register "RESERVED_CD4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F0#) =>
      -- AEB General Configuration Area Register "RESERVED_CD8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cd8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F1#) =>
      -- AEB General Configuration Area Register "RESERVED_CDC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cdc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F2#) =>
      -- AEB General Configuration Area Register "RESERVED_CE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F3#) =>
      -- AEB General Configuration Area Register "RESERVED_CE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F4#) =>
      -- AEB General Configuration Area Register "RESERVED_CE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ce8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F5#) =>
      -- AEB General Configuration Area Register "RESERVED_CEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F6#) =>
      -- AEB General Configuration Area Register "RESERVED_CF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F7#) =>
      -- AEB General Configuration Area Register "RESERVED_CF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F8#) =>
      -- AEB General Configuration Area Register "RESERVED_CF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cf8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3F9#) =>
      -- AEB General Configuration Area Register "RESERVED_CFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_cfc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FA#) =>
      -- AEB General Configuration Area Register "RESERVED_D00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FB#) =>
      -- AEB General Configuration Area Register "RESERVED_D04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FC#) =>
      -- AEB General Configuration Area Register "RESERVED_D08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FD#) =>
      -- AEB General Configuration Area Register "RESERVED_D0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FE#) =>
      -- AEB General Configuration Area Register "RESERVED_D10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#3FF#) =>
      -- AEB General Configuration Area Register "RESERVED_D14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#400#) =>
      -- AEB General Configuration Area Register "RESERVED_D18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#401#) =>
      -- AEB General Configuration Area Register "RESERVED_D1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#402#) =>
      -- AEB General Configuration Area Register "RESERVED_D20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#403#) =>
      -- AEB General Configuration Area Register "RESERVED_D24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#404#) =>
      -- AEB General Configuration Area Register "RESERVED_D28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#405#) =>
      -- AEB General Configuration Area Register "RESERVED_D2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#406#) =>
      -- AEB General Configuration Area Register "RESERVED_D30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#407#) =>
      -- AEB General Configuration Area Register "RESERVED_D34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#408#) =>
      -- AEB General Configuration Area Register "RESERVED_D38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#409#) =>
      -- AEB General Configuration Area Register "RESERVED_D3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40A#) =>
      -- AEB General Configuration Area Register "RESERVED_D40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40B#) =>
      -- AEB General Configuration Area Register "RESERVED_D44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40C#) =>
      -- AEB General Configuration Area Register "RESERVED_D48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40D#) =>
      -- AEB General Configuration Area Register "RESERVED_D4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40E#) =>
      -- AEB General Configuration Area Register "RESERVED_D50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#40F#) =>
      -- AEB General Configuration Area Register "RESERVED_D54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#410#) =>
      -- AEB General Configuration Area Register "RESERVED_D58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#411#) =>
      -- AEB General Configuration Area Register "RESERVED_D5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#412#) =>
      -- AEB General Configuration Area Register "RESERVED_D60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#413#) =>
      -- AEB General Configuration Area Register "RESERVED_D64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#414#) =>
      -- AEB General Configuration Area Register "RESERVED_D68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#415#) =>
      -- AEB General Configuration Area Register "RESERVED_D6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#416#) =>
      -- AEB General Configuration Area Register "RESERVED_D70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#417#) =>
      -- AEB General Configuration Area Register "RESERVED_D74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#418#) =>
      -- AEB General Configuration Area Register "RESERVED_D78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#419#) =>
      -- AEB General Configuration Area Register "RESERVED_D7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41A#) =>
      -- AEB General Configuration Area Register "RESERVED_D80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41B#) =>
      -- AEB General Configuration Area Register "RESERVED_D84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41C#) =>
      -- AEB General Configuration Area Register "RESERVED_D88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41D#) =>
      -- AEB General Configuration Area Register "RESERVED_D8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41E#) =>
      -- AEB General Configuration Area Register "RESERVED_D90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#41F#) =>
      -- AEB General Configuration Area Register "RESERVED_D94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#420#) =>
      -- AEB General Configuration Area Register "RESERVED_D98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#421#) =>
      -- AEB General Configuration Area Register "RESERVED_D9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_d9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#422#) =>
      -- AEB General Configuration Area Register "RESERVED_DA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#423#) =>
      -- AEB General Configuration Area Register "RESERVED_DA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#424#) =>
      -- AEB General Configuration Area Register "RESERVED_DA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_da8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#425#) =>
      -- AEB General Configuration Area Register "RESERVED_DAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#426#) =>
      -- AEB General Configuration Area Register "RESERVED_DB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#427#) =>
      -- AEB General Configuration Area Register "RESERVED_DB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#428#) =>
      -- AEB General Configuration Area Register "RESERVED_DB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_db8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#429#) =>
      -- AEB General Configuration Area Register "RESERVED_DBC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dbc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42A#) =>
      -- AEB General Configuration Area Register "RESERVED_DC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42B#) =>
      -- AEB General Configuration Area Register "RESERVED_DC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42C#) =>
      -- AEB General Configuration Area Register "RESERVED_DC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dc8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42D#) =>
      -- AEB General Configuration Area Register "RESERVED_DCC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dcc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42E#) =>
      -- AEB General Configuration Area Register "RESERVED_DD0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#42F#) =>
      -- AEB General Configuration Area Register "RESERVED_DD4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#430#) =>
      -- AEB General Configuration Area Register "RESERVED_DD8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dd8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#431#) =>
      -- AEB General Configuration Area Register "RESERVED_DDC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ddc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#432#) =>
      -- AEB General Configuration Area Register "RESERVED_DE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#433#) =>
      -- AEB General Configuration Area Register "RESERVED_DE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#434#) =>
      -- AEB General Configuration Area Register "RESERVED_DE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_de8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#435#) =>
      -- AEB General Configuration Area Register "RESERVED_DEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#436#) =>
      -- AEB General Configuration Area Register "RESERVED_DF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#437#) =>
      -- AEB General Configuration Area Register "RESERVED_DF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#438#) =>
      -- AEB General Configuration Area Register "RESERVED_DF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_df8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#439#) =>
      -- AEB General Configuration Area Register "RESERVED_DFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_dfc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43A#) =>
      -- AEB General Configuration Area Register "RESERVED_E00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43B#) =>
      -- AEB General Configuration Area Register "RESERVED_E04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43C#) =>
      -- AEB General Configuration Area Register "RESERVED_E08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43D#) =>
      -- AEB General Configuration Area Register "RESERVED_E0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43E#) =>
      -- AEB General Configuration Area Register "RESERVED_E10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#43F#) =>
      -- AEB General Configuration Area Register "RESERVED_E14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#440#) =>
      -- AEB General Configuration Area Register "RESERVED_E18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#441#) =>
      -- AEB General Configuration Area Register "RESERVED_E1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#442#) =>
      -- AEB General Configuration Area Register "RESERVED_E20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#443#) =>
      -- AEB General Configuration Area Register "RESERVED_E24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#444#) =>
      -- AEB General Configuration Area Register "RESERVED_E28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#445#) =>
      -- AEB General Configuration Area Register "RESERVED_E2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#446#) =>
      -- AEB General Configuration Area Register "RESERVED_E30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#447#) =>
      -- AEB General Configuration Area Register "RESERVED_E34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#448#) =>
      -- AEB General Configuration Area Register "RESERVED_E38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#449#) =>
      -- AEB General Configuration Area Register "RESERVED_E3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44A#) =>
      -- AEB General Configuration Area Register "RESERVED_E40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44B#) =>
      -- AEB General Configuration Area Register "RESERVED_E44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44C#) =>
      -- AEB General Configuration Area Register "RESERVED_E48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44D#) =>
      -- AEB General Configuration Area Register "RESERVED_E4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44E#) =>
      -- AEB General Configuration Area Register "RESERVED_E50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#44F#) =>
      -- AEB General Configuration Area Register "RESERVED_E54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#450#) =>
      -- AEB General Configuration Area Register "RESERVED_E58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#451#) =>
      -- AEB General Configuration Area Register "RESERVED_E5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#452#) =>
      -- AEB General Configuration Area Register "RESERVED_E60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#453#) =>
      -- AEB General Configuration Area Register "RESERVED_E64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#454#) =>
      -- AEB General Configuration Area Register "RESERVED_E68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#455#) =>
      -- AEB General Configuration Area Register "RESERVED_E6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#456#) =>
      -- AEB General Configuration Area Register "RESERVED_E70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#457#) =>
      -- AEB General Configuration Area Register "RESERVED_E74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#458#) =>
      -- AEB General Configuration Area Register "RESERVED_E78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#459#) =>
      -- AEB General Configuration Area Register "RESERVED_E7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45A#) =>
      -- AEB General Configuration Area Register "RESERVED_E80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45B#) =>
      -- AEB General Configuration Area Register "RESERVED_E84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45C#) =>
      -- AEB General Configuration Area Register "RESERVED_E88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45D#) =>
      -- AEB General Configuration Area Register "RESERVED_E8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45E#) =>
      -- AEB General Configuration Area Register "RESERVED_E90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#45F#) =>
      -- AEB General Configuration Area Register "RESERVED_E94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#460#) =>
      -- AEB General Configuration Area Register "RESERVED_E98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#461#) =>
      -- AEB General Configuration Area Register "RESERVED_E9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_e9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#462#) =>
      -- AEB General Configuration Area Register "RESERVED_EA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#463#) =>
      -- AEB General Configuration Area Register "RESERVED_EA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#464#) =>
      -- AEB General Configuration Area Register "RESERVED_EA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ea8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#465#) =>
      -- AEB General Configuration Area Register "RESERVED_EAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#466#) =>
      -- AEB General Configuration Area Register "RESERVED_EB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#467#) =>
      -- AEB General Configuration Area Register "RESERVED_EB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#468#) =>
      -- AEB General Configuration Area Register "RESERVED_EB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eb8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#469#) =>
      -- AEB General Configuration Area Register "RESERVED_EBC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ebc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46A#) =>
      -- AEB General Configuration Area Register "RESERVED_EC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46B#) =>
      -- AEB General Configuration Area Register "RESERVED_EC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46C#) =>
      -- AEB General Configuration Area Register "RESERVED_EC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ec8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46D#) =>
      -- AEB General Configuration Area Register "RESERVED_ECC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ecc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46E#) =>
      -- AEB General Configuration Area Register "RESERVED_ED0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#46F#) =>
      -- AEB General Configuration Area Register "RESERVED_ED4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#470#) =>
      -- AEB General Configuration Area Register "RESERVED_ED8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ed8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#471#) =>
      -- AEB General Configuration Area Register "RESERVED_EDC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_edc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#472#) =>
      -- AEB General Configuration Area Register "RESERVED_EE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#473#) =>
      -- AEB General Configuration Area Register "RESERVED_EE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#474#) =>
      -- AEB General Configuration Area Register "RESERVED_EE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ee8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#475#) =>
      -- AEB General Configuration Area Register "RESERVED_EEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_eec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#476#) =>
      -- AEB General Configuration Area Register "RESERVED_EF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#477#) =>
      -- AEB General Configuration Area Register "RESERVED_EF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#478#) =>
      -- AEB General Configuration Area Register "RESERVED_EF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ef8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#479#) =>
      -- AEB General Configuration Area Register "RESERVED_EFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_efc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47A#) =>
      -- AEB General Configuration Area Register "RESERVED_F00" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f00.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47B#) =>
      -- AEB General Configuration Area Register "RESERVED_F04" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f04.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47C#) =>
      -- AEB General Configuration Area Register "RESERVED_F08" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f08.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47D#) =>
      -- AEB General Configuration Area Register "RESERVED_F0C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f0c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47E#) =>
      -- AEB General Configuration Area Register "RESERVED_F10" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f10.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#47F#) =>
      -- AEB General Configuration Area Register "RESERVED_F14" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f14.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#480#) =>
      -- AEB General Configuration Area Register "RESERVED_F18" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f18.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#481#) =>
      -- AEB General Configuration Area Register "RESERVED_F1C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f1c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#482#) =>
      -- AEB General Configuration Area Register "RESERVED_F20" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f20.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#483#) =>
      -- AEB General Configuration Area Register "RESERVED_F24" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f24.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#484#) =>
      -- AEB General Configuration Area Register "RESERVED_F28" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f28.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#485#) =>
      -- AEB General Configuration Area Register "RESERVED_F2C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f2c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#486#) =>
      -- AEB General Configuration Area Register "RESERVED_F30" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f30.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#487#) =>
      -- AEB General Configuration Area Register "RESERVED_F34" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f34.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#488#) =>
      -- AEB General Configuration Area Register "RESERVED_F38" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f38.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#489#) =>
      -- AEB General Configuration Area Register "RESERVED_F3C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f3c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48A#) =>
      -- AEB General Configuration Area Register "RESERVED_F40" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f40.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48B#) =>
      -- AEB General Configuration Area Register "RESERVED_F44" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f44.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48C#) =>
      -- AEB General Configuration Area Register "RESERVED_F48" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f48.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48D#) =>
      -- AEB General Configuration Area Register "RESERVED_F4C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f4c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48E#) =>
      -- AEB General Configuration Area Register "RESERVED_F50" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f50.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#48F#) =>
      -- AEB General Configuration Area Register "RESERVED_F54" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f54.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#490#) =>
      -- AEB General Configuration Area Register "RESERVED_F58" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f58.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#491#) =>
      -- AEB General Configuration Area Register "RESERVED_F5C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f5c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#492#) =>
      -- AEB General Configuration Area Register "RESERVED_F60" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f60.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#493#) =>
      -- AEB General Configuration Area Register "RESERVED_F64" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f64.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#494#) =>
      -- AEB General Configuration Area Register "RESERVED_F68" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f68.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#495#) =>
      -- AEB General Configuration Area Register "RESERVED_F6C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f6c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#496#) =>
      -- AEB General Configuration Area Register "RESERVED_F70" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f70.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#497#) =>
      -- AEB General Configuration Area Register "RESERVED_F74" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f74.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#498#) =>
      -- AEB General Configuration Area Register "RESERVED_F78" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f78.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#499#) =>
      -- AEB General Configuration Area Register "RESERVED_F7C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f7c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49A#) =>
      -- AEB General Configuration Area Register "RESERVED_F80" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f80.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49B#) =>
      -- AEB General Configuration Area Register "RESERVED_F84" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f84.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49C#) =>
      -- AEB General Configuration Area Register "RESERVED_F88" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f88.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49D#) =>
      -- AEB General Configuration Area Register "RESERVED_F8C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f8c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49E#) =>
      -- AEB General Configuration Area Register "RESERVED_F90" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f90.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#49F#) =>
      -- AEB General Configuration Area Register "RESERVED_F94" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f94.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A0#) =>
      -- AEB General Configuration Area Register "RESERVED_F98" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f98.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A1#) =>
      -- AEB General Configuration Area Register "RESERVED_F9C" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_f9c.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A2#) =>
      -- AEB General Configuration Area Register "RESERVED_FA0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A3#) =>
      -- AEB General Configuration Area Register "RESERVED_FA4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A4#) =>
      -- AEB General Configuration Area Register "RESERVED_FA8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fa8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A5#) =>
      -- AEB General Configuration Area Register "RESERVED_FAC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fac.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A6#) =>
      -- AEB General Configuration Area Register "RESERVED_FB0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A7#) =>
      -- AEB General Configuration Area Register "RESERVED_FB4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A8#) =>
      -- AEB General Configuration Area Register "RESERVED_FB8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fb8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4A9#) =>
      -- AEB General Configuration Area Register "RESERVED_FBC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fbc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AA#) =>
      -- AEB General Configuration Area Register "RESERVED_FC0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AB#) =>
      -- AEB General Configuration Area Register "RESERVED_FC4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AC#) =>
      -- AEB General Configuration Area Register "RESERVED_FC8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fc8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AD#) =>
      -- AEB General Configuration Area Register "RESERVED_FCC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fcc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AE#) =>
      -- AEB General Configuration Area Register "RESERVED_FD0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4AF#) =>
      -- AEB General Configuration Area Register "RESERVED_FD4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B0#) =>
      -- AEB General Configuration Area Register "RESERVED_FD8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fd8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B1#) =>
      -- AEB General Configuration Area Register "RESERVED_FDC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fdc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B2#) =>
      -- AEB General Configuration Area Register "RESERVED_FE0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B3#) =>
      -- AEB General Configuration Area Register "RESERVED_FE4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B4#) =>
      -- AEB General Configuration Area Register "RESERVED_FE8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fe8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B5#) =>
      -- AEB General Configuration Area Register "RESERVED_FEC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_fec.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B6#) =>
      -- AEB General Configuration Area Register "RESERVED_FF0" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff0.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B7#) =>
      -- AEB General Configuration Area Register "RESERVED_FF4" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff4.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B8#) =>
      -- AEB General Configuration Area Register "RESERVED_FF8" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ff8.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4B9#) =>
      -- AEB General Configuration Area Register "RESERVED_FFC" : "RESERVED" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_gen_cfg_reserved_ffc.reserved(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4BA#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "AEB_STATUS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.aeb_status <= avalon_mm_rmap_i.writedata(3 downto 0);
    end if;

  when (16#4BB#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "VASP2_CFG_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.vasp2_cfg_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4BC#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "VASP1_CFG_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.vasp1_cfg_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4BD#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "DAC_CFG_WR_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.dac_cfg_wr_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4BE#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_RD_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_rd_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4BF#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_WR_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_wr_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C0#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_DAT_RD_RUN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_dat_rd_run <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C1#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_ERROR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_error <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C2#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC2_LU" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc2_lu <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C3#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC1_LU" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc1_lu <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C4#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_DAT_RD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_dat_rd <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C5#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_RD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_rd <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C6#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC_CFG_WR" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc_cfg_wr <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C7#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC2_BUSY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc2_busy <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C8#) =>
      -- AEB Housekeeping Area Register "AEB_STATUS" : "ADC1_BUSY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_aeb_status.adc1_busy <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4C9#) =>
      -- AEB Housekeeping Area Register "TIMESTAMP_1" : "TIMESTAMP_DWORD_1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_1.timestamp_dword_1(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_1.timestamp_dword_1(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_1.timestamp_dword_1(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_1.timestamp_dword_1(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4CA#) =>
      -- AEB Housekeeping Area Register "TIMESTAMP_2" : "TIMESTAMP_DWORD_0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_2.timestamp_dword_0(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_2.timestamp_dword_0(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_2.timestamp_dword_0(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_hk_timestamp_2.timestamp_dword_0(31 downto 24) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#4CB#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4CC#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4CD#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4CE#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4CF#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_L" : "ADC_CHX_DATA_T_VASP_L" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.adc_chx_data_t_vasp_l(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.adc_chx_data_t_vasp_l(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_l.adc_chx_data_t_vasp_l(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4D0#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D1#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D2#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D3#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4D4#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_VASP_R" : "ADC_CHX_DATA_T_VASP_R" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.adc_chx_data_t_vasp_r(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.adc_chx_data_t_vasp_r(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_vasp_r.adc_chx_data_t_vasp_r(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4D5#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D6#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D7#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4D8#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4D9#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_BIAS_P" : "ADC_CHX_DATA_T_BIAS_P" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.adc_chx_data_t_bias_p(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.adc_chx_data_t_bias_p(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_bias_p.adc_chx_data_t_bias_p(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4DA#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4DB#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4DC#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4DD#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4DE#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_HK_P" : "ADC_CHX_DATA_T_HK_P" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.adc_chx_data_t_hk_p(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.adc_chx_data_t_hk_p(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_hk_p.adc_chx_data_t_hk_p(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4DF#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E0#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E1#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E2#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4E3#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_1_P" : "ADC_CHX_DATA_T_TOU_1_P" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.adc_chx_data_t_tou_1_p(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.adc_chx_data_t_tou_1_p(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_1_p.adc_chx_data_t_tou_1_p(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4E4#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E5#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E6#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4E7#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4E8#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_TOU_2_P" : "ADC_CHX_DATA_T_TOU_2_P" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.adc_chx_data_t_tou_2_p(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.adc_chx_data_t_tou_2_p(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_tou_2_p.adc_chx_data_t_tou_2_p(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4E9#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4EA#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4EB#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4EC#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4ED#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODE" : "ADC_CHX_DATA_HK_VODE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.adc_chx_data_hk_vode(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.adc_chx_data_hk_vode(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vode.adc_chx_data_hk_vode(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4EE#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4EF#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F0#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F1#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4F2#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VODF" : "ADC_CHX_DATA_HK_VODF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.adc_chx_data_hk_vodf(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.adc_chx_data_hk_vodf(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vodf.adc_chx_data_hk_vodf(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4F3#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F4#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F5#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F6#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4F7#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VRD" : "ADC_CHX_DATA_HK_VRD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.adc_chx_data_hk_vrd(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.adc_chx_data_hk_vrd(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vrd.adc_chx_data_hk_vrd(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4F8#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4F9#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4FA#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4FB#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#4FC#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_VOG" : "ADC_CHX_DATA_HK_VOG" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.adc_chx_data_hk_vog(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.adc_chx_data_hk_vog(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_vog.adc_chx_data_hk_vog(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#4FD#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4FE#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#4FF#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#500#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#501#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_CCD" : "ADC_CHX_DATA_T_CCD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.adc_chx_data_t_ccd(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.adc_chx_data_t_ccd(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ccd.adc_chx_data_t_ccd(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#502#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#503#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#504#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#505#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#506#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF1K_MEA" : "ADC_CHX_DATA_T_REF1K_MEA" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.adc_chx_data_t_ref1k_mea(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.adc_chx_data_t_ref1k_mea(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref1k_mea.adc_chx_data_t_ref1k_mea(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#507#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#508#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#509#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#50A#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#50B#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_T_REF649R_MEA" : "ADC_CHX_DATA_T_REF649R_MEA" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.adc_chx_data_t_ref649r_mea(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.adc_chx_data_t_ref649r_mea(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_t_ref649r_mea.adc_chx_data_t_ref649r_mea(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#50C#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#50D#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#50E#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#50F#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#510#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_N5V" : "ADC_CHX_DATA_HK_ANA_N5V" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.adc_chx_data_hk_ana_n5v(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.adc_chx_data_hk_ana_n5v(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_n5v.adc_chx_data_hk_ana_n5v(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#511#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#512#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#513#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#514#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#515#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_S_REF" : "ADC_CHX_DATA_S_REF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.adc_chx_data_s_ref(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.adc_chx_data_s_ref(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_s_ref.adc_chx_data_s_ref(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#516#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#517#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#518#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#519#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#51A#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CCD_P31V" : "ADC_CHX_DATA_HK_CCD_P31V" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.adc_chx_data_hk_ccd_p31v(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.adc_chx_data_hk_ccd_p31v(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ccd_p31v.adc_chx_data_hk_ccd_p31v(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#51B#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#51C#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#51D#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#51E#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#51F#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_CLK_P15V" : "ADC_CHX_DATA_HK_CLK_P15V" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.adc_chx_data_hk_clk_p15v(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.adc_chx_data_hk_clk_p15v(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_clk_p15v.adc_chx_data_hk_clk_p15v(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#520#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#521#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#522#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#523#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#524#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P5V" : "ADC_CHX_DATA_HK_ANA_P5V" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.adc_chx_data_hk_ana_p5v(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.adc_chx_data_hk_ana_p5v(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p5v.adc_chx_data_hk_ana_p5v(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#525#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#526#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#527#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#528#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#529#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_ANA_P3V3" : "ADC_CHX_DATA_HK_ANA_P3V3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.adc_chx_data_hk_ana_p3v3(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.adc_chx_data_hk_ana_p3v3(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_ana_p3v3.adc_chx_data_hk_ana_p3v3(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#52A#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#52B#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#52C#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#52D#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;

  when (16#52E#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_HK_DIG_P3V3" : "ADC_CHX_DATA_HK_DIG_P3V3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.adc_chx_data_hk_dig_p3v3(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.adc_chx_data_hk_dig_p3v3(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_hk_dig_p3v3.adc_chx_data_hk_dig_p3v3(23 downto 16) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;

  when (16#52F#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "NEW" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.new_data <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#530#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "OVF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.ovf <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#531#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "SUPPLY" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.supply <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#532#) =>
      -- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "CHID" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.chid <= avalon_mm_rmap_i.writedata(4 downto 0);
    end if;
      -- AEB Housekeeping Area Register "ADC_RD_DATA_ADC_REF_BUF_2" : "ADC_CHX_DATA_ADC_REF_BUF_2" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_adc_rd_data_adc_ref_buf_2.adc_chx_data_adc_ref_buf_2 <= avalon_mm_rmap_i.writedata(11 downto 8);
    end if;

  when (16#533#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SPIRST" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.spirst <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#534#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "MUXMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.muxmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#535#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "BYPAS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.bypas <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#536#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "CLKENB" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.clkenb <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#537#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "CHOP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.chop <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#538#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "STAT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.stat <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#539#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "IDLMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.idlmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53A#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53B#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53C#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DLY0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.dly0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53D#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SBCS1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.sbcs1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53E#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "SBCS0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.sbcs0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#53F#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DRATE1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.drate1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#540#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DRATE0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.drate0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#541#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#542#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#543#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#544#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINP0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainp0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#545#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#546#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#547#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#548#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "AINN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.ainn0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#549#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54A#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54B#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54C#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54D#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54E#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#54F#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#550#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_1" : "DIFF0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_1.diff0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#551#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#552#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#553#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#554#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#555#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#556#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#557#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#558#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#559#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN15" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain15 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55A#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN14" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain14 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55B#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN13" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain13 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55C#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN12" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain12 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55D#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN11" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain11 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55E#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN10" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain10 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#55F#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN9" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain9 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#560#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "AIN8" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ain8 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#561#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "REF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.ref <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#562#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "GAIN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.gain <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#563#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "TEMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.temp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#564#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "VCC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.vcc <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#565#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "OFFSET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.offset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#566#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#567#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#568#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#569#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56A#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56B#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56C#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56D#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_2" : "CIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_2.cio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56E#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#56F#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#570#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#571#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#572#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#573#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#574#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#575#) =>
      -- AEB Housekeeping Area Register "ADC1_RD_CONFIG_3" : "DIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc1_rd_config_3.dio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#576#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SPIRST" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.spirst <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#577#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "MUXMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.muxmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#578#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "BYPAS" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.bypas <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#579#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "CLKENB" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.clkenb <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57A#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "CHOP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.chop <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57B#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "STAT" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.stat <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57C#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "IDLMOD" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.idlmod <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57D#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57E#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#57F#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DLY0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.dly0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#580#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SBCS1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.sbcs1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#581#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "SBCS0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.sbcs0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#582#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DRATE1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.drate1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#583#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DRATE0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.drate0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#584#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#585#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#586#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#587#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINP0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainp0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#588#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#589#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58A#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58B#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "AINN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.ainn0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58C#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58D#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58E#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#58F#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#590#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#591#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#592#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#593#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_1" : "DIFF0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_1.diff0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#594#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#595#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#596#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#597#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#598#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#599#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59A#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59B#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59C#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN15" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain15 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59D#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN14" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain14 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59E#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN13" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain13 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#59F#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN12" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain12 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A0#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN11" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain11 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A1#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN10" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain10 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A2#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN9" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain9 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A3#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "AIN8" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ain8 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A4#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "REF" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.ref <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A5#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "GAIN" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.gain <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A6#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "TEMP" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.temp <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A7#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "VCC" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.vcc <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A8#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "OFFSET" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.offset <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5A9#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AA#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AB#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AC#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AD#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AE#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5AF#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B0#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_2" : "CIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_2.cio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B1#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO7" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio7 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B2#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO6" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio6 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B3#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO5" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio5 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B4#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO4" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio4 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B5#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO3" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio3 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B6#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO2" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio2 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B7#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO1" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio1 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B8#) =>
      -- AEB Housekeeping Area Register "ADC2_RD_CONFIG_3" : "DIO0" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_adc2_rd_config_3.dio0 <= avalon_mm_rmap_i.writedata(0);
    end if;

  when (16#5B9#) =>
      -- AEB Housekeeping Area Register "VASP_RD_CONFIG" : "VASP1_READ_DATA" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_vasp_rd_config.vasp1_read_data <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Housekeeping Area Register "VASP_RD_CONFIG" : "VASP2_READ_DATA" Field
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_vasp_rd_config.vasp2_read_data <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Housekeeping Area Register "REVISION_ID_1" : "FPGA_VERSION" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_version(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_version(15 downto 8) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#5BA#) =>
      -- AEB Housekeeping Area Register "REVISION_ID_1" : "FPGA_DATE" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_date(7 downto 0) <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
    if (avalon_mm_rmap_i.byteenable(1) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_1.fpga_date(15 downto 8) <= avalon_mm_rmap_i.writedata(15 downto 8);
    end if;
      -- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_TIME_H" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_time_h(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_time_h(15 downto 8) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when (16#5BB#) =>
      -- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_TIME_M" Field
    if (avalon_mm_rmap_i.byteenable(0) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_time_m <= avalon_mm_rmap_i.writedata(7 downto 0);
    end if;
      -- AEB Housekeeping Area Register "REVISION_ID_2" : "FPGA_SVN" Field
    if (avalon_mm_rmap_i.byteenable(2) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_svn(7 downto 0) <= avalon_mm_rmap_i.writedata(23 downto 16);
    end if;
    if (avalon_mm_rmap_i.byteenable(3) = '1') then
      rmap_registers_wr_o.aeb_hk_revision_id_2.fpga_svn(15 downto 8) <= avalon_mm_rmap_i.writedata(31 downto 24);
    end if;

  when others =>
  -- No register associated to the address, do nothing
    null;

end case;

		end procedure p_avs_writedata;

		variable v_fee_write_address : std_logic_vector(31 downto 0)      := (others => '0');
		variable v_avs_write_address : t_farm_avalon_mm_rmap_ffee_aeb_address := 0;
	begin
		if (rst_i = '1') then
			fee_rmap_o.waitrequest       <= '1';
			avalon_mm_rmap_o.waitrequest <= '1';
			s_data_acquired              <= '0';
			p_ffee_aeb_reg_reset;
			v_fee_write_address          := (others => '0');
			v_avs_write_address          := 0;
		elsif (rising_edge(clk_i)) then

			fee_rmap_o.waitrequest       <= '1';
			avalon_mm_rmap_o.waitrequest <= '1';
			p_ffee_aeb_reg_trigger;
			s_data_acquired              <= '0';
			if (fee_rmap_i.write = '1') then
				v_fee_write_address    := fee_rmap_i.address;
				fee_rmap_o.waitrequest <= '0';
				s_data_acquired        <= '1';
				if (s_data_acquired = '0') then
					p_ffee_aeb_mem_wr(v_fee_write_address);
				end if;
			elsif (avalon_mm_rmap_i.write = '1') then
				v_avs_write_address          := to_integer(unsigned(avalon_mm_rmap_i.address));
				avalon_mm_rmap_o.waitrequest <= '0';
				s_data_acquired              <= '1';
				if (s_data_acquired = '0') then
					p_avs_writedata(v_avs_write_address);
				end if;
			end if;

		end if;
	end process p_farm_rmap_mem_area_ffee_aeb_write;

end architecture RTL;
