library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package rmap_tb_stimulli_cmd_pkg is

	-- RMAP Commands constants, subtypes and types --

	-- RMAP Commands length constants
	constant c_RMAP_CMD_13_LENGTH   : natural := 13;
	constant c_RMAP_CMD_16_LENGTH   : natural := 16;
	constant c_RMAP_CMD_17_LENGTH   : natural := 17;
	constant c_RMAP_CMD_18_LENGTH   : natural := 18;
	constant c_RMAP_CMD_22_LENGTH   : natural := 22;
	constant c_RMAP_CMD_26_LENGTH   : natural := 26;
	constant c_RMAP_CMD_274_LENGTH  : natural := 274;
	constant c_RMAP_CMD_278_LENGTH  : natural := 278;
	constant c_RMAP_CMD_4114_LENGTH : natural := 4114;
	constant c_RMAP_CMD_4118_LENGTH : natural := 4118;
	constant c_RMAP_CMD_MAX_LENGTH  : natural := 4200;

	-- RMAP Commands counter subtypes
	subtype t_rmap_cmd_13_cnt is natural range 0 to (c_RMAP_CMD_13_LENGTH - 1);
	subtype t_rmap_cmd_16_cnt is natural range 0 to (c_RMAP_CMD_16_LENGTH - 1);
	subtype t_rmap_cmd_17_cnt is natural range 0 to (c_RMAP_CMD_17_LENGTH - 1);
	subtype t_rmap_cmd_18_cnt is natural range 0 to (c_RMAP_CMD_18_LENGTH - 1);
	subtype t_rmap_cmd_22_cnt is natural range 0 to (c_RMAP_CMD_22_LENGTH - 1);
	subtype t_rmap_cmd_26_cnt is natural range 0 to (c_RMAP_CMD_26_LENGTH - 1);
	subtype t_rmap_cmd_274_cnt is natural range 0 to (c_RMAP_CMD_274_LENGTH - 1);
	subtype t_rmap_cmd_278_cnt is natural range 0 to (c_RMAP_CMD_278_LENGTH - 1);
	subtype t_rmap_cmd_4114_cnt is natural range 0 to (c_RMAP_CMD_4114_LENGTH - 1);
	subtype t_rmap_cmd_4118_cnt is natural range 0 to (c_RMAP_CMD_4118_LENGTH - 1);
	subtype t_rmap_cmd_max_cnt is natural range 0 to (c_RMAP_CMD_MAX_LENGTH - 1);

	-- RMAP Commands data types
	type t_rmap_cmd_13_data is array (0 to (c_RMAP_CMD_13_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_16_data is array (0 to (c_RMAP_CMD_16_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_17_data is array (0 to (c_RMAP_CMD_17_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_18_data is array (0 to (c_RMAP_CMD_18_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_22_data is array (0 to (c_RMAP_CMD_22_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_26_data is array (0 to (c_RMAP_CMD_26_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_274_data is array (0 to (c_RMAP_CMD_274_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_278_data is array (0 to (c_RMAP_CMD_278_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_4114_data is array (0 to (c_RMAP_CMD_4114_LENGTH - 1)) of std_logic_vector(11 downto 0);
	type t_rmap_cmd_4118_data is array (0 to (c_RMAP_CMD_4118_LENGTH - 1)) of std_logic_vector(11 downto 0);

	-- RMAP Commands test case constants --

	-- RMAP Commands test case enable constants --	
	constant c_RMAP_CMD_TEST_CASE_01_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_01_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_02_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_02_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_02_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_02_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_03_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_03_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_03_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_04_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_05_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_05_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_06_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_06_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_06_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_06_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_06_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_07_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_08_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_08_02_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_03_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_04_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_05_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_06_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_07_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_08_08_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_09_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_09_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_10_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_10_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_10_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_11_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_11_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_11_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_11_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_12_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_12_02_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_12_03_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_12_04_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_12_05_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_12_06_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_12_07_ENABLE : std_logic := '0';
	constant c_RMAP_CMD_TEST_CASE_13_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_13_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_13_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_13_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_13_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_13_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_13_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_14_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_15_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_16_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_17_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_18_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_19_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_20_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_21_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_22_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_23_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_24_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_25_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_14_26_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_15_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_15_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_15_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_15_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_15_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_16_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_16_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_16_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_16_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_13_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_14_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_15_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_16_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_17_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_17_18_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_13_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_14_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_15_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_16_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_17_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_18_18_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_13_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_14_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_15_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_16_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_17_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_19_18_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_01_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_02_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_03_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_04_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_05_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_06_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_07_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_08_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_09_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_10_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_11_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_12_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_13_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_14_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_15_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_16_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_17_ENABLE : std_logic := '1';
	constant c_RMAP_CMD_TEST_CASE_20_18_ENABLE : std_logic := '1';

	-- RMAP Commands test case times constants --	
	constant c_RMAP_CMD_TEST_CASE_01_01_TIME : natural := 100;
	constant c_RMAP_CMD_TEST_CASE_01_02_TIME : natural := 200;
	constant c_RMAP_CMD_TEST_CASE_01_03_TIME : natural := 300;
	constant c_RMAP_CMD_TEST_CASE_01_04_TIME : natural := 400;
	constant c_RMAP_CMD_TEST_CASE_01_05_TIME : natural := 500;
	constant c_RMAP_CMD_TEST_CASE_01_06_TIME : natural := 600;
	constant c_RMAP_CMD_TEST_CASE_01_07_TIME : natural := 700;
	constant c_RMAP_CMD_TEST_CASE_02_01_TIME : natural := 800;
	constant c_RMAP_CMD_TEST_CASE_02_02_TIME : natural := 900;
	constant c_RMAP_CMD_TEST_CASE_02_03_TIME : natural := 1000;
	constant c_RMAP_CMD_TEST_CASE_02_04_TIME : natural := 1100;
	constant c_RMAP_CMD_TEST_CASE_03_01_TIME : natural := 1200;
	constant c_RMAP_CMD_TEST_CASE_03_02_TIME : natural := 1300;
	constant c_RMAP_CMD_TEST_CASE_03_03_TIME : natural := 1400;
	constant c_RMAP_CMD_TEST_CASE_04_01_TIME : natural := 1500;
	constant c_RMAP_CMD_TEST_CASE_04_02_TIME : natural := 1600;
	constant c_RMAP_CMD_TEST_CASE_04_03_TIME : natural := 1700;
	constant c_RMAP_CMD_TEST_CASE_04_04_TIME : natural := 1800;
	constant c_RMAP_CMD_TEST_CASE_04_05_TIME : natural := 1900;
	constant c_RMAP_CMD_TEST_CASE_04_06_TIME : natural := 2000;
	constant c_RMAP_CMD_TEST_CASE_04_07_TIME : natural := 2100;
	constant c_RMAP_CMD_TEST_CASE_04_08_TIME : natural := 2200;
	constant c_RMAP_CMD_TEST_CASE_04_09_TIME : natural := 2300;
	constant c_RMAP_CMD_TEST_CASE_04_10_TIME : natural := 2400;
	constant c_RMAP_CMD_TEST_CASE_04_11_TIME : natural := 2500;
	constant c_RMAP_CMD_TEST_CASE_04_12_TIME : natural := 2600;
	constant c_RMAP_CMD_TEST_CASE_05_01_TIME : natural := 2700;
	constant c_RMAP_CMD_TEST_CASE_05_02_TIME : natural := 2800;
	constant c_RMAP_CMD_TEST_CASE_06_01_TIME : natural := 2900;
	constant c_RMAP_CMD_TEST_CASE_06_02_TIME : natural := 3000;
	constant c_RMAP_CMD_TEST_CASE_06_03_TIME : natural := 3100;
	constant c_RMAP_CMD_TEST_CASE_06_04_TIME : natural := 3200;
	constant c_RMAP_CMD_TEST_CASE_06_05_TIME : natural := 3300;
	constant c_RMAP_CMD_TEST_CASE_07_01_TIME : natural := 3400;
	constant c_RMAP_CMD_TEST_CASE_07_02_TIME : natural := 3500;
	constant c_RMAP_CMD_TEST_CASE_07_03_TIME : natural := 3600;
	constant c_RMAP_CMD_TEST_CASE_07_04_TIME : natural := 3700;
	constant c_RMAP_CMD_TEST_CASE_07_05_TIME : natural := 3800;
	constant c_RMAP_CMD_TEST_CASE_07_06_TIME : natural := 3900;
	constant c_RMAP_CMD_TEST_CASE_07_07_TIME : natural := 4000;
	constant c_RMAP_CMD_TEST_CASE_07_08_TIME : natural := 4100;
	constant c_RMAP_CMD_TEST_CASE_07_09_TIME : natural := 4200;
	constant c_RMAP_CMD_TEST_CASE_07_10_TIME : natural := 4300;
	constant c_RMAP_CMD_TEST_CASE_08_01_TIME : natural := 4400;
	constant c_RMAP_CMD_TEST_CASE_08_02_TIME : natural := 4500;
	constant c_RMAP_CMD_TEST_CASE_08_03_TIME : natural := 4600;
	constant c_RMAP_CMD_TEST_CASE_08_04_TIME : natural := 4700;
	constant c_RMAP_CMD_TEST_CASE_08_05_TIME : natural := 4800;
	constant c_RMAP_CMD_TEST_CASE_08_06_TIME : natural := 4900;
	constant c_RMAP_CMD_TEST_CASE_08_07_TIME : natural := 5000;
	constant c_RMAP_CMD_TEST_CASE_08_08_TIME : natural := 5100;
	constant c_RMAP_CMD_TEST_CASE_09_01_TIME : natural := 5200;
	constant c_RMAP_CMD_TEST_CASE_09_02_TIME : natural := 5300;
	constant c_RMAP_CMD_TEST_CASE_09_03_TIME : natural := 5400;
	constant c_RMAP_CMD_TEST_CASE_09_04_TIME : natural := 5500;
	constant c_RMAP_CMD_TEST_CASE_09_05_TIME : natural := 5600;
	constant c_RMAP_CMD_TEST_CASE_09_06_TIME : natural := 5700;
	constant c_RMAP_CMD_TEST_CASE_09_07_TIME : natural := 5800;
	constant c_RMAP_CMD_TEST_CASE_09_08_TIME : natural := 5900;
	constant c_RMAP_CMD_TEST_CASE_09_09_TIME : natural := 6000;
	constant c_RMAP_CMD_TEST_CASE_09_10_TIME : natural := 6100;
	constant c_RMAP_CMD_TEST_CASE_10_01_TIME : natural := 6200;
	constant c_RMAP_CMD_TEST_CASE_10_02_TIME : natural := 6300;
	constant c_RMAP_CMD_TEST_CASE_10_03_TIME : natural := 6400;
	constant c_RMAP_CMD_TEST_CASE_11_01_TIME : natural := 6500;
	constant c_RMAP_CMD_TEST_CASE_11_02_TIME : natural := 6600;
	constant c_RMAP_CMD_TEST_CASE_11_03_TIME : natural := 6700;
	constant c_RMAP_CMD_TEST_CASE_11_04_TIME : natural := 6800;
	constant c_RMAP_CMD_TEST_CASE_12_01_TIME : natural := 6900;
	constant c_RMAP_CMD_TEST_CASE_12_02_TIME : natural := 7000;
	constant c_RMAP_CMD_TEST_CASE_12_03_TIME : natural := 7100;
	constant c_RMAP_CMD_TEST_CASE_12_04_TIME : natural := 7200;
	constant c_RMAP_CMD_TEST_CASE_12_05_TIME : natural := 7300;
	constant c_RMAP_CMD_TEST_CASE_12_06_TIME : natural := 7400;
	constant c_RMAP_CMD_TEST_CASE_12_07_TIME : natural := 7500;
	constant c_RMAP_CMD_TEST_CASE_13_01_TIME : natural := 7600;
	constant c_RMAP_CMD_TEST_CASE_13_02_TIME : natural := 7700;
	constant c_RMAP_CMD_TEST_CASE_13_03_TIME : natural := 7800;
	constant c_RMAP_CMD_TEST_CASE_13_04_TIME : natural := 7900;
	constant c_RMAP_CMD_TEST_CASE_13_05_TIME : natural := 8000;
	constant c_RMAP_CMD_TEST_CASE_13_06_TIME : natural := 8100;
	constant c_RMAP_CMD_TEST_CASE_14_01_TIME : natural := 8200;
	constant c_RMAP_CMD_TEST_CASE_14_02_TIME : natural := 8300;
	constant c_RMAP_CMD_TEST_CASE_14_03_TIME : natural := 8400;
	constant c_RMAP_CMD_TEST_CASE_14_04_TIME : natural := 8500;
	constant c_RMAP_CMD_TEST_CASE_14_05_TIME : natural := 8600;
	constant c_RMAP_CMD_TEST_CASE_14_06_TIME : natural := 8700;
	constant c_RMAP_CMD_TEST_CASE_14_07_TIME : natural := 8800;
	constant c_RMAP_CMD_TEST_CASE_14_08_TIME : natural := 8900;
	constant c_RMAP_CMD_TEST_CASE_14_09_TIME : natural := 9000;
	constant c_RMAP_CMD_TEST_CASE_14_10_TIME : natural := 9100;
	constant c_RMAP_CMD_TEST_CASE_14_11_TIME : natural := 9200;
	constant c_RMAP_CMD_TEST_CASE_14_12_TIME : natural := 9300;
	constant c_RMAP_CMD_TEST_CASE_14_13_TIME : natural := 9400;
	constant c_RMAP_CMD_TEST_CASE_14_14_TIME : natural := 9500;
	constant c_RMAP_CMD_TEST_CASE_14_15_TIME : natural := 9600;
	constant c_RMAP_CMD_TEST_CASE_14_16_TIME : natural := 9700;
	constant c_RMAP_CMD_TEST_CASE_14_17_TIME : natural := 9800;
	constant c_RMAP_CMD_TEST_CASE_14_18_TIME : natural := 9900;
	constant c_RMAP_CMD_TEST_CASE_14_19_TIME : natural := 10000;
	constant c_RMAP_CMD_TEST_CASE_14_20_TIME : natural := 10100;
	constant c_RMAP_CMD_TEST_CASE_14_21_TIME : natural := 10200;
	constant c_RMAP_CMD_TEST_CASE_14_22_TIME : natural := 10300;
	constant c_RMAP_CMD_TEST_CASE_14_23_TIME : natural := 10400;
	constant c_RMAP_CMD_TEST_CASE_14_24_TIME : natural := 10500;
	constant c_RMAP_CMD_TEST_CASE_14_25_TIME : natural := 10600;
	constant c_RMAP_CMD_TEST_CASE_14_26_TIME : natural := 10700;
	constant c_RMAP_CMD_TEST_CASE_15_01_TIME : natural := 10800;
	constant c_RMAP_CMD_TEST_CASE_15_02_TIME : natural := 10900;
	constant c_RMAP_CMD_TEST_CASE_15_03_TIME : natural := 11000;
	constant c_RMAP_CMD_TEST_CASE_15_04_TIME : natural := 11100;
	constant c_RMAP_CMD_TEST_CASE_15_05_TIME : natural := 11200;
	constant c_RMAP_CMD_TEST_CASE_16_01_TIME : natural := 11300;
	constant c_RMAP_CMD_TEST_CASE_16_02_TIME : natural := 11400;
	constant c_RMAP_CMD_TEST_CASE_16_03_TIME : natural := 11500;
	constant c_RMAP_CMD_TEST_CASE_16_04_TIME : natural := 11600;
	constant c_RMAP_CMD_TEST_CASE_17_01_TIME : natural := 11700;
	constant c_RMAP_CMD_TEST_CASE_17_02_TIME : natural := 11800;
	constant c_RMAP_CMD_TEST_CASE_17_03_TIME : natural := 11900;
	constant c_RMAP_CMD_TEST_CASE_17_04_TIME : natural := 12000;
	constant c_RMAP_CMD_TEST_CASE_17_05_TIME : natural := 12100;
	constant c_RMAP_CMD_TEST_CASE_17_06_TIME : natural := 12200;
	constant c_RMAP_CMD_TEST_CASE_17_07_TIME : natural := 12300;
	constant c_RMAP_CMD_TEST_CASE_17_08_TIME : natural := 12400;
	constant c_RMAP_CMD_TEST_CASE_17_09_TIME : natural := 12500;
	constant c_RMAP_CMD_TEST_CASE_17_10_TIME : natural := 12600;
	constant c_RMAP_CMD_TEST_CASE_17_11_TIME : natural := 12700;
	constant c_RMAP_CMD_TEST_CASE_17_12_TIME : natural := 12800;
	constant c_RMAP_CMD_TEST_CASE_17_13_TIME : natural := 12900;
	constant c_RMAP_CMD_TEST_CASE_17_14_TIME : natural := 13000;
	constant c_RMAP_CMD_TEST_CASE_17_15_TIME : natural := 13100;
	constant c_RMAP_CMD_TEST_CASE_17_16_TIME : natural := 13200;
	constant c_RMAP_CMD_TEST_CASE_17_17_TIME : natural := 13300;
	constant c_RMAP_CMD_TEST_CASE_17_18_TIME : natural := 13400;
	constant c_RMAP_CMD_TEST_CASE_18_01_TIME : natural := 13500;
	constant c_RMAP_CMD_TEST_CASE_18_02_TIME : natural := 13600;
	constant c_RMAP_CMD_TEST_CASE_18_03_TIME : natural := 13700;
	constant c_RMAP_CMD_TEST_CASE_18_04_TIME : natural := 13800;
	constant c_RMAP_CMD_TEST_CASE_18_05_TIME : natural := 13900;
	constant c_RMAP_CMD_TEST_CASE_18_06_TIME : natural := 14000;
	constant c_RMAP_CMD_TEST_CASE_18_07_TIME : natural := 14100;
	constant c_RMAP_CMD_TEST_CASE_18_08_TIME : natural := 14200;
	constant c_RMAP_CMD_TEST_CASE_18_09_TIME : natural := 14300;
	constant c_RMAP_CMD_TEST_CASE_18_10_TIME : natural := 14400;
	constant c_RMAP_CMD_TEST_CASE_18_11_TIME : natural := 14500;
	constant c_RMAP_CMD_TEST_CASE_18_12_TIME : natural := 14600;
	constant c_RMAP_CMD_TEST_CASE_18_13_TIME : natural := 14700;
	constant c_RMAP_CMD_TEST_CASE_18_14_TIME : natural := 14800;
	constant c_RMAP_CMD_TEST_CASE_18_15_TIME : natural := 14900;
	constant c_RMAP_CMD_TEST_CASE_18_16_TIME : natural := 15000;
	constant c_RMAP_CMD_TEST_CASE_18_17_TIME : natural := 15100;
	constant c_RMAP_CMD_TEST_CASE_18_18_TIME : natural := 15200;
	constant c_RMAP_CMD_TEST_CASE_19_01_TIME : natural := 15300;
	constant c_RMAP_CMD_TEST_CASE_19_02_TIME : natural := 15400;
	constant c_RMAP_CMD_TEST_CASE_19_03_TIME : natural := 15500;
	constant c_RMAP_CMD_TEST_CASE_19_04_TIME : natural := 15600;
	constant c_RMAP_CMD_TEST_CASE_19_05_TIME : natural := 15700;
	constant c_RMAP_CMD_TEST_CASE_19_06_TIME : natural := 15800;
	constant c_RMAP_CMD_TEST_CASE_19_07_TIME : natural := 15900;
	constant c_RMAP_CMD_TEST_CASE_19_08_TIME : natural := 16000;
	constant c_RMAP_CMD_TEST_CASE_19_09_TIME : natural := 16100;
	constant c_RMAP_CMD_TEST_CASE_19_10_TIME : natural := 16200;
	constant c_RMAP_CMD_TEST_CASE_19_11_TIME : natural := 16300;
	constant c_RMAP_CMD_TEST_CASE_19_12_TIME : natural := 16400;
	constant c_RMAP_CMD_TEST_CASE_19_13_TIME : natural := 16500;
	constant c_RMAP_CMD_TEST_CASE_19_14_TIME : natural := 16600;
	constant c_RMAP_CMD_TEST_CASE_19_15_TIME : natural := 16700;
	constant c_RMAP_CMD_TEST_CASE_19_16_TIME : natural := 16800;
	constant c_RMAP_CMD_TEST_CASE_19_17_TIME : natural := 16900;
	constant c_RMAP_CMD_TEST_CASE_19_18_TIME : natural := 17000;
	constant c_RMAP_CMD_TEST_CASE_20_01_TIME : natural := 17100;
	constant c_RMAP_CMD_TEST_CASE_20_02_TIME : natural := 17200;
	constant c_RMAP_CMD_TEST_CASE_20_03_TIME : natural := 17300;
	constant c_RMAP_CMD_TEST_CASE_20_04_TIME : natural := 17400;
	constant c_RMAP_CMD_TEST_CASE_20_05_TIME : natural := 17500;
	constant c_RMAP_CMD_TEST_CASE_20_06_TIME : natural := 17600;
	constant c_RMAP_CMD_TEST_CASE_20_07_TIME : natural := 17700;
	constant c_RMAP_CMD_TEST_CASE_20_08_TIME : natural := 17800;
	constant c_RMAP_CMD_TEST_CASE_20_09_TIME : natural := 17900;
	constant c_RMAP_CMD_TEST_CASE_20_10_TIME : natural := 18000;
	constant c_RMAP_CMD_TEST_CASE_20_11_TIME : natural := 18100;
	constant c_RMAP_CMD_TEST_CASE_20_12_TIME : natural := 18200;
	constant c_RMAP_CMD_TEST_CASE_20_13_TIME : natural := 18300;
	constant c_RMAP_CMD_TEST_CASE_20_14_TIME : natural := 18400;
	constant c_RMAP_CMD_TEST_CASE_20_15_TIME : natural := 18500;
	constant c_RMAP_CMD_TEST_CASE_20_16_TIME : natural := 18600;
	constant c_RMAP_CMD_TEST_CASE_20_17_TIME : natural := 18700;
	constant c_RMAP_CMD_TEST_CASE_20_18_TIME : natural := 18800;
	constant c_RMAP_CMD_TEST_FINISH_TIME     : natural := 18900;

	-- RMAP Commands test case text constants --	
	constant c_RMAP_CMD_TEST_CASE_01_01_TEXT : string := "RMAP Test Case 1.1";
	constant c_RMAP_CMD_TEST_CASE_01_02_TEXT : string := "RMAP Test Case 1.2";
	constant c_RMAP_CMD_TEST_CASE_01_03_TEXT : string := "RMAP Test Case 1.3";
	constant c_RMAP_CMD_TEST_CASE_01_04_TEXT : string := "RMAP Test Case 1.4";
	constant c_RMAP_CMD_TEST_CASE_01_05_TEXT : string := "RMAP Test Case 1.5";
	constant c_RMAP_CMD_TEST_CASE_01_06_TEXT : string := "RMAP Test Case 1.6";
	constant c_RMAP_CMD_TEST_CASE_01_07_TEXT : string := "RMAP Test Case 1.7";
	constant c_RMAP_CMD_TEST_CASE_02_01_TEXT : string := "RMAP Test Case 2.1";
	constant c_RMAP_CMD_TEST_CASE_02_02_TEXT : string := "RMAP Test Case 2.2";
	constant c_RMAP_CMD_TEST_CASE_02_03_TEXT : string := "RMAP Test Case 2.3";
	constant c_RMAP_CMD_TEST_CASE_02_04_TEXT : string := "RMAP Test Case 2.4";
	constant c_RMAP_CMD_TEST_CASE_03_01_TEXT : string := "RMAP Test Case 3.1";
	constant c_RMAP_CMD_TEST_CASE_03_02_TEXT : string := "RMAP Test Case 3.2";
	constant c_RMAP_CMD_TEST_CASE_03_03_TEXT : string := "RMAP Test Case 3.3";
	constant c_RMAP_CMD_TEST_CASE_04_01_TEXT : string := "RMAP Test Case 4.1";
	constant c_RMAP_CMD_TEST_CASE_04_02_TEXT : string := "RMAP Test Case 4.2";
	constant c_RMAP_CMD_TEST_CASE_04_03_TEXT : string := "RMAP Test Case 4.3";
	constant c_RMAP_CMD_TEST_CASE_04_04_TEXT : string := "RMAP Test Case 4.4";
	constant c_RMAP_CMD_TEST_CASE_04_05_TEXT : string := "RMAP Test Case 4.5";
	constant c_RMAP_CMD_TEST_CASE_04_06_TEXT : string := "RMAP Test Case 4.6";
	constant c_RMAP_CMD_TEST_CASE_04_07_TEXT : string := "RMAP Test Case 4.7";
	constant c_RMAP_CMD_TEST_CASE_04_08_TEXT : string := "RMAP Test Case 4.8";
	constant c_RMAP_CMD_TEST_CASE_04_09_TEXT : string := "RMAP Test Case 4.9";
	constant c_RMAP_CMD_TEST_CASE_04_10_TEXT : string := "RMAP Test Case 4.10";
	constant c_RMAP_CMD_TEST_CASE_04_11_TEXT : string := "RMAP Test Case 4.11";
	constant c_RMAP_CMD_TEST_CASE_04_12_TEXT : string := "RMAP Test Case 4.12";
	constant c_RMAP_CMD_TEST_CASE_05_01_TEXT : string := "RMAP Test Case 5.1";
	constant c_RMAP_CMD_TEST_CASE_05_02_TEXT : string := "RMAP Test Case 5.2";
	constant c_RMAP_CMD_TEST_CASE_06_01_TEXT : string := "RMAP Test Case 6.1";
	constant c_RMAP_CMD_TEST_CASE_06_02_TEXT : string := "RMAP Test Case 6.2";
	constant c_RMAP_CMD_TEST_CASE_06_03_TEXT : string := "RMAP Test Case 6.3";
	constant c_RMAP_CMD_TEST_CASE_06_04_TEXT : string := "RMAP Test Case 6.4";
	constant c_RMAP_CMD_TEST_CASE_06_05_TEXT : string := "RMAP Test Case 6.5";
	constant c_RMAP_CMD_TEST_CASE_07_01_TEXT : string := "RMAP Test Case 7.1";
	constant c_RMAP_CMD_TEST_CASE_07_02_TEXT : string := "RMAP Test Case 7.2";
	constant c_RMAP_CMD_TEST_CASE_07_03_TEXT : string := "RMAP Test Case 7.3";
	constant c_RMAP_CMD_TEST_CASE_07_04_TEXT : string := "RMAP Test Case 7.4";
	constant c_RMAP_CMD_TEST_CASE_07_05_TEXT : string := "RMAP Test Case 7.5";
	constant c_RMAP_CMD_TEST_CASE_07_06_TEXT : string := "RMAP Test Case 7.6";
	constant c_RMAP_CMD_TEST_CASE_07_07_TEXT : string := "RMAP Test Case 7.7";
	constant c_RMAP_CMD_TEST_CASE_07_08_TEXT : string := "RMAP Test Case 7.8";
	constant c_RMAP_CMD_TEST_CASE_07_09_TEXT : string := "RMAP Test Case 7.9";
	constant c_RMAP_CMD_TEST_CASE_07_10_TEXT : string := "RMAP Test Case 7.10";
	constant c_RMAP_CMD_TEST_CASE_08_01_TEXT : string := "RMAP Test Case 8.1";
	constant c_RMAP_CMD_TEST_CASE_08_02_TEXT : string := "RMAP Test Case 8.2";
	constant c_RMAP_CMD_TEST_CASE_08_03_TEXT : string := "RMAP Test Case 8.3";
	constant c_RMAP_CMD_TEST_CASE_08_04_TEXT : string := "RMAP Test Case 8.4";
	constant c_RMAP_CMD_TEST_CASE_08_05_TEXT : string := "RMAP Test Case 8.5";
	constant c_RMAP_CMD_TEST_CASE_08_06_TEXT : string := "RMAP Test Case 8.6";
	constant c_RMAP_CMD_TEST_CASE_08_07_TEXT : string := "RMAP Test Case 8.7";
	constant c_RMAP_CMD_TEST_CASE_08_08_TEXT : string := "RMAP Test Case 8.8";
	constant c_RMAP_CMD_TEST_CASE_09_01_TEXT : string := "RMAP Test Case 9.1";
	constant c_RMAP_CMD_TEST_CASE_09_02_TEXT : string := "RMAP Test Case 9.2";
	constant c_RMAP_CMD_TEST_CASE_09_03_TEXT : string := "RMAP Test Case 9.3";
	constant c_RMAP_CMD_TEST_CASE_09_04_TEXT : string := "RMAP Test Case 9.4";
	constant c_RMAP_CMD_TEST_CASE_09_05_TEXT : string := "RMAP Test Case 9.5";
	constant c_RMAP_CMD_TEST_CASE_09_06_TEXT : string := "RMAP Test Case 9.6";
	constant c_RMAP_CMD_TEST_CASE_09_07_TEXT : string := "RMAP Test Case 9.7";
	constant c_RMAP_CMD_TEST_CASE_09_08_TEXT : string := "RMAP Test Case 9.8";
	constant c_RMAP_CMD_TEST_CASE_09_09_TEXT : string := "RMAP Test Case 9.9";
	constant c_RMAP_CMD_TEST_CASE_09_10_TEXT : string := "RMAP Test Case 9.10";
	constant c_RMAP_CMD_TEST_CASE_10_01_TEXT : string := "RMAP Test Case 10.1";
	constant c_RMAP_CMD_TEST_CASE_10_02_TEXT : string := "RMAP Test Case 10.2";
	constant c_RMAP_CMD_TEST_CASE_10_03_TEXT : string := "RMAP Test Case 10.3";
	constant c_RMAP_CMD_TEST_CASE_11_01_TEXT : string := "RMAP Test Case 11.1";
	constant c_RMAP_CMD_TEST_CASE_11_02_TEXT : string := "RMAP Test Case 11.2";
	constant c_RMAP_CMD_TEST_CASE_11_03_TEXT : string := "RMAP Test Case 11.3";
	constant c_RMAP_CMD_TEST_CASE_11_04_TEXT : string := "RMAP Test Case 11.4";
	constant c_RMAP_CMD_TEST_CASE_12_01_TEXT : string := "RMAP Test Case 12.1";
	constant c_RMAP_CMD_TEST_CASE_12_02_TEXT : string := "RMAP Test Case 12.2";
	constant c_RMAP_CMD_TEST_CASE_12_03_TEXT : string := "RMAP Test Case 12.3";
	constant c_RMAP_CMD_TEST_CASE_12_04_TEXT : string := "RMAP Test Case 12.4";
	constant c_RMAP_CMD_TEST_CASE_12_05_TEXT : string := "RMAP Test Case 12.5";
	constant c_RMAP_CMD_TEST_CASE_12_06_TEXT : string := "RMAP Test Case 12.6";
	constant c_RMAP_CMD_TEST_CASE_12_07_TEXT : string := "RMAP Test Case 12.7";
	constant c_RMAP_CMD_TEST_CASE_13_01_TEXT : string := "RMAP Test Case 13.1";
	constant c_RMAP_CMD_TEST_CASE_13_02_TEXT : string := "RMAP Test Case 13.2";
	constant c_RMAP_CMD_TEST_CASE_13_03_TEXT : string := "RMAP Test Case 13.3";
	constant c_RMAP_CMD_TEST_CASE_13_04_TEXT : string := "RMAP Test Case 13.4";
	constant c_RMAP_CMD_TEST_CASE_13_05_TEXT : string := "RMAP Test Case 13.5";
	constant c_RMAP_CMD_TEST_CASE_13_06_TEXT : string := "RMAP Test Case 13.6";
	constant c_RMAP_CMD_TEST_CASE_14_01_TEXT : string := "RMAP Test Case 14.1";
	constant c_RMAP_CMD_TEST_CASE_14_02_TEXT : string := "RMAP Test Case 14.2";
	constant c_RMAP_CMD_TEST_CASE_14_03_TEXT : string := "RMAP Test Case 14.3";
	constant c_RMAP_CMD_TEST_CASE_14_04_TEXT : string := "RMAP Test Case 14.4";
	constant c_RMAP_CMD_TEST_CASE_14_05_TEXT : string := "RMAP Test Case 14.5";
	constant c_RMAP_CMD_TEST_CASE_14_06_TEXT : string := "RMAP Test Case 14.6";
	constant c_RMAP_CMD_TEST_CASE_14_07_TEXT : string := "RMAP Test Case 14.7";
	constant c_RMAP_CMD_TEST_CASE_14_08_TEXT : string := "RMAP Test Case 14.8";
	constant c_RMAP_CMD_TEST_CASE_14_09_TEXT : string := "RMAP Test Case 14.9";
	constant c_RMAP_CMD_TEST_CASE_14_10_TEXT : string := "RMAP Test Case 14.10";
	constant c_RMAP_CMD_TEST_CASE_14_11_TEXT : string := "RMAP Test Case 14.11";
	constant c_RMAP_CMD_TEST_CASE_14_12_TEXT : string := "RMAP Test Case 14.12";
	constant c_RMAP_CMD_TEST_CASE_14_13_TEXT : string := "RMAP Test Case 14.13";
	constant c_RMAP_CMD_TEST_CASE_14_14_TEXT : string := "RMAP Test Case 14.14";
	constant c_RMAP_CMD_TEST_CASE_14_15_TEXT : string := "RMAP Test Case 14.15";
	constant c_RMAP_CMD_TEST_CASE_14_16_TEXT : string := "RMAP Test Case 14.16";
	constant c_RMAP_CMD_TEST_CASE_14_17_TEXT : string := "RMAP Test Case 14.17";
	constant c_RMAP_CMD_TEST_CASE_14_18_TEXT : string := "RMAP Test Case 14.18";
	constant c_RMAP_CMD_TEST_CASE_14_19_TEXT : string := "RMAP Test Case 14.19";
	constant c_RMAP_CMD_TEST_CASE_14_20_TEXT : string := "RMAP Test Case 14.20";
	constant c_RMAP_CMD_TEST_CASE_14_21_TEXT : string := "RMAP Test Case 14.21";
	constant c_RMAP_CMD_TEST_CASE_14_22_TEXT : string := "RMAP Test Case 14.22";
	constant c_RMAP_CMD_TEST_CASE_14_23_TEXT : string := "RMAP Test Case 14.23";
	constant c_RMAP_CMD_TEST_CASE_14_24_TEXT : string := "RMAP Test Case 14.24";
	constant c_RMAP_CMD_TEST_CASE_14_25_TEXT : string := "RMAP Test Case 14.25";
	constant c_RMAP_CMD_TEST_CASE_14_26_TEXT : string := "RMAP Test Case 14.26";
	constant c_RMAP_CMD_TEST_CASE_15_01_TEXT : string := "RMAP Test Case 15.1";
	constant c_RMAP_CMD_TEST_CASE_15_02_TEXT : string := "RMAP Test Case 15.2";
	constant c_RMAP_CMD_TEST_CASE_15_03_TEXT : string := "RMAP Test Case 15.3";
	constant c_RMAP_CMD_TEST_CASE_15_04_TEXT : string := "RMAP Test Case 15.4";
	constant c_RMAP_CMD_TEST_CASE_15_05_TEXT : string := "RMAP Test Case 15.5";
	constant c_RMAP_CMD_TEST_CASE_16_01_TEXT : string := "RMAP Test Case 16.1";
	constant c_RMAP_CMD_TEST_CASE_16_02_TEXT : string := "RMAP Test Case 16.2";
	constant c_RMAP_CMD_TEST_CASE_16_03_TEXT : string := "RMAP Test Case 16.3";
	constant c_RMAP_CMD_TEST_CASE_16_04_TEXT : string := "RMAP Test Case 16.4";
	constant c_RMAP_CMD_TEST_CASE_17_01_TEXT : string := "RMAP Test Case 17.1";
	constant c_RMAP_CMD_TEST_CASE_17_02_TEXT : string := "RMAP Test Case 17.2";
	constant c_RMAP_CMD_TEST_CASE_17_03_TEXT : string := "RMAP Test Case 17.3";
	constant c_RMAP_CMD_TEST_CASE_17_04_TEXT : string := "RMAP Test Case 17.4";
	constant c_RMAP_CMD_TEST_CASE_17_05_TEXT : string := "RMAP Test Case 17.5";
	constant c_RMAP_CMD_TEST_CASE_17_06_TEXT : string := "RMAP Test Case 17.6";
	constant c_RMAP_CMD_TEST_CASE_17_07_TEXT : string := "RMAP Test Case 17.7";
	constant c_RMAP_CMD_TEST_CASE_17_08_TEXT : string := "RMAP Test Case 17.8";
	constant c_RMAP_CMD_TEST_CASE_17_09_TEXT : string := "RMAP Test Case 17.9";
	constant c_RMAP_CMD_TEST_CASE_17_10_TEXT : string := "RMAP Test Case 17.10";
	constant c_RMAP_CMD_TEST_CASE_17_11_TEXT : string := "RMAP Test Case 17.11";
	constant c_RMAP_CMD_TEST_CASE_17_12_TEXT : string := "RMAP Test Case 17.12";
	constant c_RMAP_CMD_TEST_CASE_17_13_TEXT : string := "RMAP Test Case 17.13";
	constant c_RMAP_CMD_TEST_CASE_17_14_TEXT : string := "RMAP Test Case 17.14";
	constant c_RMAP_CMD_TEST_CASE_17_15_TEXT : string := "RMAP Test Case 17.15";
	constant c_RMAP_CMD_TEST_CASE_17_16_TEXT : string := "RMAP Test Case 17.16";
	constant c_RMAP_CMD_TEST_CASE_17_17_TEXT : string := "RMAP Test Case 17.17";
	constant c_RMAP_CMD_TEST_CASE_17_18_TEXT : string := "RMAP Test Case 17.18";
	constant c_RMAP_CMD_TEST_CASE_18_01_TEXT : string := "RMAP Test Case 18.1";
	constant c_RMAP_CMD_TEST_CASE_18_02_TEXT : string := "RMAP Test Case 18.2";
	constant c_RMAP_CMD_TEST_CASE_18_03_TEXT : string := "RMAP Test Case 18.3";
	constant c_RMAP_CMD_TEST_CASE_18_04_TEXT : string := "RMAP Test Case 18.4";
	constant c_RMAP_CMD_TEST_CASE_18_05_TEXT : string := "RMAP Test Case 18.5";
	constant c_RMAP_CMD_TEST_CASE_18_06_TEXT : string := "RMAP Test Case 18.6";
	constant c_RMAP_CMD_TEST_CASE_18_07_TEXT : string := "RMAP Test Case 18.7";
	constant c_RMAP_CMD_TEST_CASE_18_08_TEXT : string := "RMAP Test Case 18.8";
	constant c_RMAP_CMD_TEST_CASE_18_09_TEXT : string := "RMAP Test Case 18.9";
	constant c_RMAP_CMD_TEST_CASE_18_10_TEXT : string := "RMAP Test Case 18.10";
	constant c_RMAP_CMD_TEST_CASE_18_11_TEXT : string := "RMAP Test Case 18.11";
	constant c_RMAP_CMD_TEST_CASE_18_12_TEXT : string := "RMAP Test Case 18.12";
	constant c_RMAP_CMD_TEST_CASE_18_13_TEXT : string := "RMAP Test Case 18.13";
	constant c_RMAP_CMD_TEST_CASE_18_14_TEXT : string := "RMAP Test Case 18.14";
	constant c_RMAP_CMD_TEST_CASE_18_15_TEXT : string := "RMAP Test Case 18.15";
	constant c_RMAP_CMD_TEST_CASE_18_16_TEXT : string := "RMAP Test Case 18.16";
	constant c_RMAP_CMD_TEST_CASE_18_17_TEXT : string := "RMAP Test Case 18.17";
	constant c_RMAP_CMD_TEST_CASE_18_18_TEXT : string := "RMAP Test Case 18.18";
	constant c_RMAP_CMD_TEST_CASE_19_01_TEXT : string := "RMAP Test Case 19.1";
	constant c_RMAP_CMD_TEST_CASE_19_02_TEXT : string := "RMAP Test Case 19.2";
	constant c_RMAP_CMD_TEST_CASE_19_03_TEXT : string := "RMAP Test Case 19.3";
	constant c_RMAP_CMD_TEST_CASE_19_04_TEXT : string := "RMAP Test Case 19.4";
	constant c_RMAP_CMD_TEST_CASE_19_05_TEXT : string := "RMAP Test Case 19.5";
	constant c_RMAP_CMD_TEST_CASE_19_06_TEXT : string := "RMAP Test Case 19.6";
	constant c_RMAP_CMD_TEST_CASE_19_07_TEXT : string := "RMAP Test Case 19.7";
	constant c_RMAP_CMD_TEST_CASE_19_08_TEXT : string := "RMAP Test Case 19.8";
	constant c_RMAP_CMD_TEST_CASE_19_09_TEXT : string := "RMAP Test Case 19.9";
	constant c_RMAP_CMD_TEST_CASE_19_10_TEXT : string := "RMAP Test Case 19.10";
	constant c_RMAP_CMD_TEST_CASE_19_11_TEXT : string := "RMAP Test Case 19.11";
	constant c_RMAP_CMD_TEST_CASE_19_12_TEXT : string := "RMAP Test Case 19.12";
	constant c_RMAP_CMD_TEST_CASE_19_13_TEXT : string := "RMAP Test Case 19.13";
	constant c_RMAP_CMD_TEST_CASE_19_14_TEXT : string := "RMAP Test Case 19.14";
	constant c_RMAP_CMD_TEST_CASE_19_15_TEXT : string := "RMAP Test Case 19.15";
	constant c_RMAP_CMD_TEST_CASE_19_16_TEXT : string := "RMAP Test Case 19.16";
	constant c_RMAP_CMD_TEST_CASE_19_17_TEXT : string := "RMAP Test Case 19.17";
	constant c_RMAP_CMD_TEST_CASE_19_18_TEXT : string := "RMAP Test Case 19.18";
	constant c_RMAP_CMD_TEST_CASE_20_01_TEXT : string := "RMAP Test Case 20.1";
	constant c_RMAP_CMD_TEST_CASE_20_02_TEXT : string := "RMAP Test Case 20.2";
	constant c_RMAP_CMD_TEST_CASE_20_03_TEXT : string := "RMAP Test Case 20.3";
	constant c_RMAP_CMD_TEST_CASE_20_04_TEXT : string := "RMAP Test Case 20.4";
	constant c_RMAP_CMD_TEST_CASE_20_05_TEXT : string := "RMAP Test Case 20.5";
	constant c_RMAP_CMD_TEST_CASE_20_06_TEXT : string := "RMAP Test Case 20.6";
	constant c_RMAP_CMD_TEST_CASE_20_07_TEXT : string := "RMAP Test Case 20.7";
	constant c_RMAP_CMD_TEST_CASE_20_08_TEXT : string := "RMAP Test Case 20.8";
	constant c_RMAP_CMD_TEST_CASE_20_09_TEXT : string := "RMAP Test Case 20.9";
	constant c_RMAP_CMD_TEST_CASE_20_10_TEXT : string := "RMAP Test Case 20.10";
	constant c_RMAP_CMD_TEST_CASE_20_11_TEXT : string := "RMAP Test Case 20.11";
	constant c_RMAP_CMD_TEST_CASE_20_12_TEXT : string := "RMAP Test Case 20.12";
	constant c_RMAP_CMD_TEST_CASE_20_13_TEXT : string := "RMAP Test Case 20.13";
	constant c_RMAP_CMD_TEST_CASE_20_14_TEXT : string := "RMAP Test Case 20.14";
	constant c_RMAP_CMD_TEST_CASE_20_15_TEXT : string := "RMAP Test Case 20.15";
	constant c_RMAP_CMD_TEST_CASE_20_16_TEXT : string := "RMAP Test Case 20.16";
	constant c_RMAP_CMD_TEST_CASE_20_17_TEXT : string := "RMAP Test Case 20.17";
	constant c_RMAP_CMD_TEST_CASE_20_18_TEXT : string := "RMAP Test Case 20.18";

	-- RMAP Commands test case data constants

	-- Test Case 1.1 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Correct Protocol ID = 0x01 RMAP Protocol 
	constant c_RMAP_CMD_TEST_CASE_01_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 1.2 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0x02 CCSDS Packet Encapsulation Protocol 
	constant c_RMAP_CMD_TEST_CASE_01_02_DATA : t_rmap_cmd_17_data   := (x"051", x"002", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0E3", x"100");
	-- Test Case 1.3 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0x00 Extended Protocol Identifier 
	constant c_RMAP_CMD_TEST_CASE_01_03_DATA : t_rmap_cmd_17_data   := (x"051", x"000", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"014", x"100");
	-- Test Case 1.4 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0x03 
	constant c_RMAP_CMD_TEST_CASE_01_04_DATA : t_rmap_cmd_17_data   := (x"051", x"003", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"078", x"100");
	-- Test Case 1.5 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0x11 
	constant c_RMAP_CMD_TEST_CASE_01_05_DATA : t_rmap_cmd_17_data   := (x"051", x"011", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"033", x"100");
	-- Test Case 1.6 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0xEE GOES-R Reliable Data Delivery Protocol 
	constant c_RMAP_CMD_TEST_CASE_01_06_DATA : t_rmap_cmd_17_data   := (x"051", x"0EE", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"03F", x"100");
	-- Test Case 1.7 (PLATO-DLR-PL-ICD-0007 4.5.1.9): Wrong protocol ID = 0xEF Serial Transfer Universal Protocol 
	constant c_RMAP_CMD_TEST_CASE_01_07_DATA : t_rmap_cmd_17_data   := (x"051", x"0EF", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0A4", x"100");
	-- Test Case 2.1 (PLATO-DLR-PL-ICD-0007 4.1): Correct reply address length
	constant c_RMAP_CMD_TEST_CASE_02_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 2.2 (PLATO-DLR-PL-ICD-0007 4.1): Reply Address length check = 1
	constant c_RMAP_CMD_TEST_CASE_02_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04D", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"000", x"100");
	-- Test Case 2.3 (PLATO-DLR-PL-ICD-0007 4.1): Reply Address length check = 2
	constant c_RMAP_CMD_TEST_CASE_02_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04E", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"050", x"100");
	-- Test Case 2.4 (PLATO-DLR-PL-ICD-0007 4.1): Reply Address length check = 3
	constant c_RMAP_CMD_TEST_CASE_02_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04F", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0DF", x"100");
	-- Test Case 3.1 (PLATO-DLR-PL-ICD-0007 4.5.1.5): Valid read packet with EOP
	constant c_RMAP_CMD_TEST_CASE_03_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 3.2 (PLATO-DLR-PL-ICD-0007 4.5.1.5): Invalid read packet with EEP
	constant c_RMAP_CMD_TEST_CASE_03_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0FB", x"101");
	-- Test Case 3.3 (PLATO-DLR-PL-ICD-0007 4.5.1.5): Invalid write packet with EEP
	constant c_RMAP_CMD_TEST_CASE_03_03_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"008", x"05A", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"101");
	-- Test Case 4.1 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Valid command code 0x4C
	constant c_RMAP_CMD_TEST_CASE_04_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 4.2 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Valid command code 0x6C
	constant c_RMAP_CMD_TEST_CASE_04_02_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"07F", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 4.3 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 0x6C to critical memory 0x00000014
	constant c_RMAP_CMD_TEST_CASE_04_03_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"0D3", x"000", x"000", x"000", x"006", x"0E4", x"100");
	-- Test Case 4.4 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 0x6C to housekeeping memory 0x00001000
	constant c_RMAP_CMD_TEST_CASE_04_04_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"010", x"000", x"000", x"000", x"004", x"0F1", x"000", x"000", x"000", x"006", x"0E4", x"100");
	-- Test Case 4.5 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Valid command code 0x7C
	constant c_RMAP_CMD_TEST_CASE_04_05_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"006", x"000", x"000", x"000", x"006", x"0E4", x"100");
	-- Test Case 4.6 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 0x7C to housekeeping memory 0x00001000
	constant c_RMAP_CMD_TEST_CASE_04_06_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"000", x"010", x"000", x"000", x"000", x"004", x"094", x"006", x"000", x"000", x"000", x"0AA", x"100");
	-- Test Case 4.7 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 0
	constant c_RMAP_CMD_TEST_CASE_04_07_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"040", x"0D1", x"050", x"000", x"007", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0E6", x"100");
	-- Test Case 4.8 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 1
	constant c_RMAP_CMD_TEST_CASE_04_08_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"044", x"0D1", x"050", x"000", x"008", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0FC", x"100");
	-- Test Case 4.9 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 4
	constant c_RMAP_CMD_TEST_CASE_04_09_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"050", x"0D1", x"050", x"000", x"009", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"092", x"100");
	-- Test Case 4.10 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 5
	constant c_RMAP_CMD_TEST_CASE_04_10_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"054", x"0D1", x"050", x"000", x"00A", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"099", x"100");
	-- Test Case 4.11 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 6
	constant c_RMAP_CMD_TEST_CASE_04_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"058", x"0D1", x"050", x"000", x"00B", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"034", x"100");
	-- Test Case 4.12 (PLATO-DLR-PL-ICD-0007 4.5.1.10): Invalid command code 7
	constant c_RMAP_CMD_TEST_CASE_04_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"05C", x"0D1", x"050", x"000", x"00C", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 5.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): No data characters in read command
	constant c_RMAP_CMD_TEST_CASE_05_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 5.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Data characters in read command
	constant c_RMAP_CMD_TEST_CASE_05_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"008", x"0F2", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 6.1 (PLATO-DLR-PL-ICD-0007 4.5.1.7): Valid Key = 0xD1
	constant c_RMAP_CMD_TEST_CASE_06_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 6.2 (PLATO-DLR-PL-ICD-0007 4.5.1.7): Invalid Key = 0xD0
	constant c_RMAP_CMD_TEST_CASE_06_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D0", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0A9", x"100");
	-- Test Case 6.3 (PLATO-DLR-PL-ICD-0007 4.5.1.7): Invalid Key = 0xD2
	constant c_RMAP_CMD_TEST_CASE_06_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D2", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"021", x"100");
	-- Test Case 6.4 (PLATO-DLR-PL-ICD-0007 4.5.1.7): Invalid Key = 0x00
	constant c_RMAP_CMD_TEST_CASE_06_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"000", x"050", x"000", x"004", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0C1", x"100");
	-- Test Case 6.5 (PLATO-DLR-PL-ICD-0007 4.5.1.7): Invalid Key = 0xFF
	constant c_RMAP_CMD_TEST_CASE_06_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0FF", x"050", x"000", x"005", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"00F", x"100");
	-- Test Case 7.1 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Valid logical target address = 0x51
	constant c_RMAP_CMD_TEST_CASE_07_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 7.2 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x00
	constant c_RMAP_CMD_TEST_CASE_07_02_DATA : t_rmap_cmd_17_data   := (x"000", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"000", x"100");
	-- Test Case 7.3 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0xFF
	constant c_RMAP_CMD_TEST_CASE_07_03_DATA : t_rmap_cmd_17_data   := (x"0FF", x"001", x"04C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"025", x"100");
	-- Test Case 7.4 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x61
	constant c_RMAP_CMD_TEST_CASE_07_04_DATA : t_rmap_cmd_17_data   := (x"061", x"001", x"04C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"085", x"100");
	-- Test Case 7.5 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x41
	constant c_RMAP_CMD_TEST_CASE_07_05_DATA : t_rmap_cmd_17_data   := (x"041", x"001", x"04C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0F2", x"100");
	-- Test Case 7.6 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0xFE
	constant c_RMAP_CMD_TEST_CASE_07_06_DATA : t_rmap_cmd_17_data   := (x"0FE", x"001", x"04C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"039", x"100");
	-- Test Case 7.7 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x11
	constant c_RMAP_CMD_TEST_CASE_07_07_DATA : t_rmap_cmd_17_data   := (x"011", x"001", x"04C", x"0D1", x"050", x"000", x"007", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0D1", x"100");
	-- Test Case 7.8 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x99
	constant c_RMAP_CMD_TEST_CASE_07_08_DATA : t_rmap_cmd_17_data   := (x"099", x"001", x"04C", x"0D1", x"050", x"000", x"008", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"09F", x"100");
	-- Test Case 7.9 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x50
	constant c_RMAP_CMD_TEST_CASE_07_09_DATA : t_rmap_cmd_17_data   := (x"050", x"001", x"04C", x"0D1", x"050", x"000", x"009", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0AE", x"100");
	-- Test Case 7.10 (PLATO-DLR-PL-ICD-0007 4.5.1.8): Invalid logical target address = 0x52
	constant c_RMAP_CMD_TEST_CASE_07_10_DATA : t_rmap_cmd_17_data   := (x"052", x"001", x"04C", x"0D1", x"050", x"000", x"00A", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"01B", x"100");
	-- Test Case 8.1 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from valid address
	constant c_RMAP_CMD_TEST_CASE_08_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 8.2 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused address 0x00090000
	constant c_RMAP_CMD_TEST_CASE_08_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"009", x"000", x"000", x"000", x"000", x"004", x"0B5", x"100");
	-- Test Case 8.3 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused address 0x10000000
	constant c_RMAP_CMD_TEST_CASE_08_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"003", x"000", x"010", x"000", x"000", x"000", x"000", x"000", x"004", x"080", x"100");
	-- Test Case 8.4 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused DEB address 0x00008000
	constant c_RMAP_CMD_TEST_CASE_08_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"080", x"000", x"000", x"000", x"004", x"055", x"100");
	-- Test Case 8.5 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused AEB1 address 0x00018000
	constant c_RMAP_CMD_TEST_CASE_08_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"001", x"080", x"000", x"000", x"000", x"004", x"04E", x"100");
	-- Test Case 8.6 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused AEB2 address 0x00028000
	constant c_RMAP_CMD_TEST_CASE_08_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"002", x"080", x"000", x"000", x"000", x"004", x"063", x"100");
	-- Test Case 8.7 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused AEB3 address 0x00048000
	constant c_RMAP_CMD_TEST_CASE_08_07_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"007", x"000", x"000", x"004", x"080", x"000", x"000", x"000", x"004", x"0FD", x"100");
	-- Test Case 8.8 (PLATO-DLR-PL-ICD-0007 4.5.1.3): Read from unused AEB4 address 0x00088000
	constant c_RMAP_CMD_TEST_CASE_08_08_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"008", x"000", x"000", x"008", x"080", x"000", x"000", x"000", x"004", x"03D", x"100");
	-- Test Case 9.1 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Valid header
	constant c_RMAP_CMD_TEST_CASE_09_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 9.2 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Header CRC Error - overwrite header crc to 0x00
	constant c_RMAP_CMD_TEST_CASE_09_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"000", x"100");
	-- Test Case 9.3 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Header CRC Error - overwrite header crc to 0xFF
	constant c_RMAP_CMD_TEST_CASE_09_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0FF", x"100");
	-- Test Case 9.4 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Incomplete header - remove protocol ID
	constant c_RMAP_CMD_TEST_CASE_09_04_DATA : t_rmap_cmd_16_data   := (x"051", x"04C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"013", x"100");
	-- Test Case 9.5 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Incomplete header - remove key
	constant c_RMAP_CMD_TEST_CASE_09_05_DATA : t_rmap_cmd_16_data   := (x"051", x"001", x"04C", x"050", x"000", x"005", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"03F", x"100");
	-- Test Case 9.6 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Incomplete header - remove first address byte (MSB)
	constant c_RMAP_CMD_TEST_CASE_09_06_DATA : t_rmap_cmd_16_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"04B", x"100");
	-- Test Case 9.7 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Incomplete header - remove all address bytes
	constant c_RMAP_CMD_TEST_CASE_09_07_DATA : t_rmap_cmd_13_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"007", x"000", x"000", x"000", x"004", x"067", x"100");
	-- Test Case 9.8 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Invalid header - Unused packet type = 0
	constant c_RMAP_CMD_TEST_CASE_09_08_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"00C", x"0D1", x"050", x"000", x"008", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"0F6", x"100");
	-- Test Case 9.9 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Invalid header - Unused packet type = 2
	constant c_RMAP_CMD_TEST_CASE_09_09_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"0CC", x"0D1", x"050", x"000", x"009", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"007", x"100");
	-- Test Case 9.10 (PLATO-DLR-PL-ICD-0007 4.5.1.4): Invalid header - Unused packet type = 3
	constant c_RMAP_CMD_TEST_CASE_09_10_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"0CC", x"0D1", x"050", x"000", x"00A", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"073", x"100");
	-- Test Case 10.1 (PLATO-DLR-PL-ICD-0007 4.5.1.6): Valid Data CRC
	constant c_RMAP_CMD_TEST_CASE_10_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"00B", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 10.2 (PLATO-DLR-PL-ICD-0007 4.5.1.6): Invalid Data CRC 0x00
	constant c_RMAP_CMD_TEST_CASE_10_02_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"07F", x"000", x"000", x"000", x"0EE", x"000", x"100");
	-- Test Case 10.3 (PLATO-DLR-PL-ICD-0007 4.5.1.6): Invalid Data CRC 0xFF
	constant c_RMAP_CMD_TEST_CASE_10_03_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"053", x"000", x"000", x"000", x"0EE", x"0FF", x"100");
	-- Test Case 11.1 (PLATO-DLR-PL-ICD-0007 4.5.1.1): Write to valid address 0x00000130
	constant c_RMAP_CMD_TEST_CASE_11_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"00B", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 11.2 (PLATO-DLR-PL-ICD-0007 4.5.1.1): Write 8 Bytes across memory border starting at address 0x000000FC
	constant c_RMAP_CMD_TEST_CASE_11_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"0FC", x"000", x"000", x"008", x"06B", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 11.3 (PLATO-DLR-PL-ICD-0007 4.5.1.1): Write 8 Bytes across memory border starting at address 0x00000FFC
	constant c_RMAP_CMD_TEST_CASE_11_03_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"00F", x"0FC", x"000", x"000", x"008", x"0EA", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 11.4 (PLATO-DLR-PL-ICD-0007 4.5.1.1): Write 8 Bytes across memory border starting at address 0x00001FFC
	constant c_RMAP_CMD_TEST_CASE_11_04_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"01F", x"0FC", x"000", x"000", x"008", x"0B6", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 12.1 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to valid address 0x00000130
	constant c_RMAP_CMD_TEST_CASE_12_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"00B", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.2 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused address 0x10000000
	constant c_RMAP_CMD_TEST_CASE_12_02_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"002", x"000", x"010", x"000", x"000", x"000", x"000", x"000", x"004", x"0D6", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.3 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused DEB address 0x00008000
	constant c_RMAP_CMD_TEST_CASE_12_03_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"080", x"000", x"000", x"000", x"004", x"0EB", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.4 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused AEB1 address 0x00018000
	constant c_RMAP_CMD_TEST_CASE_12_04_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"001", x"080", x"000", x"000", x"000", x"004", x"018", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.5 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused AEB2 address 0x00028000
	constant c_RMAP_CMD_TEST_CASE_12_05_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"002", x"080", x"000", x"000", x"000", x"004", x"06D", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.6 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused AEB3 address 0x00048000
	constant c_RMAP_CMD_TEST_CASE_12_06_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"004", x"080", x"000", x"000", x"000", x"004", x"0AB", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 12.7 (PLATO-DLR-PL-ICD-0007 4.5.1.2): Write to unused AEB4 address 0x00088000
	constant c_RMAP_CMD_TEST_CASE_12_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"007", x"000", x"000", x"001", x"080", x"000", x"000", x"000", x"004", x"06C", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 13.1 (PLATO-DLR-PL-ICD-0007 4.5.1.11): Correct amount of data
	constant c_RMAP_CMD_TEST_CASE_13_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"00B", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 13.2 (PLATO-DLR-PL-ICD-0007 4.5.1.11): Less data than expected (expected 8 Bytes; provided 4 Bytes)
	constant c_RMAP_CMD_TEST_CASE_13_02_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"008", x"076", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 13.3 (PLATO-DLR-PL-ICD-0007 4.5.1.11): Less data than expected (expected 260 Bytes; provided 4 Bytes)
	constant c_RMAP_CMD_TEST_CASE_13_03_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"001", x"030", x"000", x"001", x"004", x"03E", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 13.4 (PLATO-DLR-PL-ICD-0007 4.5.1.11): Less data than expected (expected 16777212 Bytes; provided 4 Bytes)
	constant c_RMAP_CMD_TEST_CASE_13_04_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"001", x"030", x"0FF", x"0FF", x"0FC", x"012", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 13.5 (PLATO-DLR-PL-ICD-0007 4.5.1.11): More data than expected (expected 4 Bytes; provided 8 Bytes)
	constant c_RMAP_CMD_TEST_CASE_13_05_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"0BB", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 13.6 (PLATO-DLR-PL-ICD-0007 4.5.1.11): More data than expected (expected 0 Bytes; provided 4 Bytes)
	constant c_RMAP_CMD_TEST_CASE_13_06_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"000", x"0C8", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 14.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 bytes to DEB critical configuration are (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"0B6", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 14.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 8 Bytes to DEB critical configuration area (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"008", x"0CB", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 14.3 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to DEB critical configuration area (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_03_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"000", x"0E9", x"000", x"100");
	-- Test Case 14.4 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 4 Bytes from DEB critical configuration area (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"06D", x"100");
	-- Test Case 14.5 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 8 Bytes from DEB critical configuration area (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"008", x"048", x"100");
	-- Test Case 14.6 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 0 Bytes from DEB critical configuration area (0x00000014)
	constant c_RMAP_CMD_TEST_CASE_14_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"006", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"000", x"032", x"100");
	-- Test Case 14.7 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"007", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"0E3", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 14.8 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 256 Bytes to DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_08_DATA : t_rmap_cmd_274_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"008", x"000", x"000", x"000", x"001", x"030", x"000", x"001", x"000", x"0EC", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"0A9", x"100");
	-- Test Case 14.9 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 260 Bytes to DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_09_DATA : t_rmap_cmd_278_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"009", x"000", x"000", x"000", x"001", x"030", x"000", x"001", x"004", x"0C7", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"018", x"100");
	-- Test Case 14.10 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_10_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"00A", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"000", x"0D9", x"000", x"100");
	-- Test Case 14.11 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"00B", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"088", x"100");
	-- Test Case 14.12 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"00C", x"000", x"000", x"000", x"001", x"030", x"000", x"001", x"000", x"026", x"100");
	-- Test Case 14.13 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_13_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"00D", x"000", x"000", x"000", x"001", x"030", x"000", x"001", x"004", x"00D", x"100");
	-- Test Case 14.14 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from DEB general configuration area (0x00000130)
	constant c_RMAP_CMD_TEST_CASE_14_14_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"00E", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"000", x"013", x"100");
	-- Test Case 14.15 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from DEB housekeeping area (0x00001000)
	constant c_RMAP_CMD_TEST_CASE_14_15_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"00F", x"000", x"000", x"000", x"010", x"000", x"000", x"000", x"004", x"05E", x"100");
	-- Test Case 14.16 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from DEB housekeeping area (0x00001000)
	constant c_RMAP_CMD_TEST_CASE_14_16_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"010", x"000", x"000", x"000", x"010", x"000", x"000", x"001", x"000", x"0D2", x"100");
	-- Test Case 14.17 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from DEB housekeeping area (0x00001000)
	constant c_RMAP_CMD_TEST_CASE_14_17_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"011", x"000", x"000", x"000", x"010", x"000", x"000", x"001", x"004", x"0F9", x"100");
	-- Test Case 14.18 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from DEB housekeeping area (0x00001000)
	constant c_RMAP_CMD_TEST_CASE_14_18_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"012", x"000", x"000", x"000", x"010", x"000", x"000", x"000", x"000", x"0E7", x"100");
	-- Test Case 14.19 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_19_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"013", x"000", x"000", x"000", x"020", x"000", x"000", x"000", x"004", x"0DF", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 14.20 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4096 Bytes to DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_20_DATA : t_rmap_cmd_4114_data := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"014", x"000", x"000", x"000", x"020", x"000", x"000", x"010", x"000", x"009", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"08D", x"100");
	-- Test Case 14.21 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4100 Bytes to DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_21_DATA : t_rmap_cmd_4118_data := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"015", x"000", x"000", x"000", x"020", x"000", x"000", x"010", x"004", x"022", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"071", x"100");
	-- Test Case 14.22 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_22_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"016", x"000", x"000", x"000", x"020", x"000", x"000", x"000", x"000", x"044", x"000", x"100");
	-- Test Case 14.23 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_23_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"017", x"000", x"000", x"000", x"020", x"000", x"000", x"000", x"004", x"015", x"100");
	-- Test Case 14.24 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4096 Bytes from DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_24_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"018", x"000", x"000", x"000", x"020", x"000", x"000", x"010", x"000", x"062", x"100");
	-- Test Case 14.25 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4100 Bytes from DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_25_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"019", x"000", x"000", x"000", x"020", x"000", x"000", x"010", x"004", x"049", x"100");
	-- Test Case 14.26 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from DEB windowing area (0x00002000)
	constant c_RMAP_CMD_TEST_CASE_14_26_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"01A", x"000", x"000", x"000", x"020", x"000", x"000", x"000", x"000", x"02F", x"100");
	-- Test Case 15.1 (PLATO-DLR-PL-ICD-0007 4.5.1.13): Valid 4-Byte aligned data length field
	constant c_RMAP_CMD_TEST_CASE_15_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"004", x"08F", x"100");
	-- Test Case 15.2 (PLATO-DLR-PL-ICD-0007 4.5.1.13): Invalid aligned data length field: 3 Bytes
	constant c_RMAP_CMD_TEST_CASE_15_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"003", x"08E", x"100");
	-- Test Case 15.3 (PLATO-DLR-PL-ICD-0007 4.5.1.13): Invalid aligned data length field: 5 Bytes
	constant c_RMAP_CMD_TEST_CASE_15_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"005", x"046", x"100");
	-- Test Case 15.4 (PLATO-DLR-PL-ICD-0007 4.5.1.13): Invalid aligned data length field: 6 Bytes
	constant c_RMAP_CMD_TEST_CASE_15_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"006", x"0F0", x"100");
	-- Test Case 15.5 (PLATO-DLR-PL-ICD-0007 4.5.1.13): Invalid aligned data length field: 14 Bytes
	constant c_RMAP_CMD_TEST_CASE_15_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"005", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"00E", x"02C", x"100");
	-- Test Case 16.1 (PLATO-DLR-PL-ICD-0007 4.1 / 4.5.1.10): Valid read with incrementing address
	constant c_RMAP_CMD_TEST_CASE_16_01_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"001", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"0F1", x"100");
	-- Test Case 16.2 (PLATO-DLR-PL-ICD-0007 4.1 / 4.5.1.10): Invalid read without incrementing address
	constant c_RMAP_CMD_TEST_CASE_16_02_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"048", x"0D1", x"050", x"000", x"002", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"0FA", x"100");
	-- Test Case 16.3 (PLATO-DLR-PL-ICD-0007 4.1 / 4.5.1.10): Invalid verified write without incrementing address
	constant c_RMAP_CMD_TEST_CASE_16_03_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"078", x"0D1", x"050", x"000", x"003", x"000", x"000", x"000", x"000", x"014", x"000", x"000", x"004", x"091", x"100");
	-- Test Case 16.4 (PLATO-DLR-PL-ICD-0007 4.1 / 4.5.1.10): Invalid unverified write without incrementing address
	constant c_RMAP_CMD_TEST_CASE_16_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"068", x"0D1", x"050", x"000", x"004", x"000", x"000", x"000", x"001", x"030", x"000", x"000", x"004", x"0E8", x"100");
	-- Test Case 17.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 bytes to AEB1 critical configuration are (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"01B", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"004", x"0FB", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 17.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 8 Bytes to AEB1 critical configuration area (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"01C", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"008", x"036", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 17.3 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB1 critical configuration area (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_03_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"01D", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"000", x"014", x"000", x"100");
	-- Test Case 17.4 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 4 Bytes from AEB1 critical configuration area (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"01E", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"004", x"020", x"100");
	-- Test Case 17.5 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 8 Bytes from AEB1 critical configuration area (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"01F", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"008", x"005", x"100");
	-- Test Case 17.6 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 0 Bytes from AEB1 critical configuration area (0x00010014)
	constant c_RMAP_CMD_TEST_CASE_17_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"020", x"000", x"000", x"001", x"000", x"014", x"000", x"000", x"000", x"02A", x"100");
	-- Test Case 17.7 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"021", x"000", x"000", x"001", x"001", x"030", x"000", x"000", x"004", x"0FB", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 17.8 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 256 Bytes to AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_08_DATA : t_rmap_cmd_274_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"022", x"000", x"000", x"001", x"001", x"030", x"000", x"001", x"000", x"0E5", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"0A9", x"100");
	-- Test Case 17.9 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 260 Bytes to AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_09_DATA : t_rmap_cmd_278_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"023", x"000", x"000", x"001", x"001", x"030", x"000", x"001", x"004", x"0CE", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"018", x"100");
	-- Test Case 17.10 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_10_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"024", x"000", x"000", x"001", x"001", x"030", x"000", x"000", x"000", x"060", x"000", x"100");
	-- Test Case 17.11 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"025", x"000", x"000", x"001", x"001", x"030", x"000", x"000", x"004", x"031", x"100");
	-- Test Case 17.12 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"026", x"000", x"000", x"001", x"001", x"030", x"000", x"001", x"000", x"02F", x"100");
	-- Test Case 17.13 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_13_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"027", x"000", x"000", x"001", x"001", x"030", x"000", x"001", x"004", x"004", x"100");
	-- Test Case 17.14 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB1 general configuration area (0x00010130)
	constant c_RMAP_CMD_TEST_CASE_17_14_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"028", x"000", x"000", x"001", x"001", x"030", x"000", x"000", x"000", x"00B", x"100");
	-- Test Case 17.15 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB1 housekeeping area (0x00011000)
	constant c_RMAP_CMD_TEST_CASE_17_15_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"029", x"000", x"000", x"001", x"010", x"000", x"000", x"000", x"004", x"046", x"100");
	-- Test Case 17.16 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB1 housekeeping area (0x00011000)
	constant c_RMAP_CMD_TEST_CASE_17_16_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"02A", x"000", x"000", x"001", x"010", x"000", x"000", x"001", x"000", x"058", x"100");
	-- Test Case 17.17 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB1 housekeeping area (0x00011000)
	constant c_RMAP_CMD_TEST_CASE_17_17_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"02B", x"000", x"000", x"001", x"010", x"000", x"000", x"001", x"004", x"073", x"100");
	-- Test Case 17.18 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB1 housekeeping area (0x00011000)
	constant c_RMAP_CMD_TEST_CASE_17_18_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"02C", x"000", x"000", x"001", x"010", x"000", x"000", x"000", x"000", x"0DD", x"100");
	-- Test Case 18.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 bytes to AEB2 critical configuration are (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"02D", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"004", x"00E", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 18.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 8 Bytes to AEB2 critical configuration area (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"02E", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"008", x"073", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 18.3 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB2 critical configuration area (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_03_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"02F", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"000", x"051", x"000", x"100");
	-- Test Case 18.4 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 4 Bytes from AEB2 critical configuration area (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"030", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"004", x"0F7", x"100");
	-- Test Case 18.5 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 8 Bytes from AEB2 critical configuration area (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"031", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"008", x"0D2", x"100");
	-- Test Case 18.6 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 0 Bytes from AEB2 critical configuration area (0x00020014)
	constant c_RMAP_CMD_TEST_CASE_18_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"032", x"000", x"000", x"002", x"000", x"014", x"000", x"000", x"000", x"0A8", x"100");
	-- Test Case 18.7 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"033", x"000", x"000", x"002", x"001", x"030", x"000", x"000", x"004", x"079", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 18.8 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 256 Bytes to AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_08_DATA : t_rmap_cmd_274_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"034", x"000", x"000", x"002", x"001", x"030", x"000", x"001", x"000", x"0D7", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"0A9", x"100");
	-- Test Case 18.9 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 260 Bytes to AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_09_DATA : t_rmap_cmd_278_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"035", x"000", x"000", x"002", x"001", x"030", x"000", x"001", x"004", x"0FC", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"018", x"100");
	-- Test Case 18.10 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_10_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"036", x"000", x"000", x"002", x"001", x"030", x"000", x"000", x"000", x"0E2", x"000", x"100");
	-- Test Case 18.11 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"037", x"000", x"000", x"002", x"001", x"030", x"000", x"000", x"004", x"0B3", x"100");
	-- Test Case 18.12 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"038", x"000", x"000", x"002", x"001", x"030", x"000", x"001", x"000", x"0BC", x"100");
	-- Test Case 18.13 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_13_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"039", x"000", x"000", x"002", x"001", x"030", x"000", x"001", x"004", x"097", x"100");
	-- Test Case 18.14 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB2 general configuration area (0x00020130)
	constant c_RMAP_CMD_TEST_CASE_18_14_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"03A", x"000", x"000", x"002", x"001", x"030", x"000", x"000", x"000", x"089", x"100");
	-- Test Case 18.15 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB2 housekeeping area (0x00021000)
	constant c_RMAP_CMD_TEST_CASE_18_15_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"03B", x"000", x"000", x"002", x"010", x"000", x"000", x"000", x"004", x"0C4", x"100");
	-- Test Case 18.16 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB2 housekeeping area (0x00021000)
	constant c_RMAP_CMD_TEST_CASE_18_16_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"03C", x"000", x"000", x"002", x"010", x"000", x"000", x"001", x"000", x"06A", x"100");
	-- Test Case 18.17 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB2 housekeeping area (0x00021000)
	constant c_RMAP_CMD_TEST_CASE_18_17_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"03D", x"000", x"000", x"002", x"010", x"000", x"000", x"001", x"004", x"041", x"100");
	-- Test Case 18.18 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB2 housekeeping area (0x00021000)
	constant c_RMAP_CMD_TEST_CASE_18_18_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"03E", x"000", x"000", x"002", x"010", x"000", x"000", x"000", x"000", x"05F", x"100");
	-- Test Case 19.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 bytes to AEB3 critical configuration are (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"03F", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"004", x"067", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 19.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 8 Bytes to AEB3 critical configuration area (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"040", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"008", x"000", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 19.3 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB3 critical configuration area (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_03_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"041", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"000", x"022", x"000", x"100");
	-- Test Case 19.4 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 4 Bytes from AEB3 critical configuration area (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"042", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"004", x"016", x"100");
	-- Test Case 19.5 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 8 Bytes from AEB3 critical configuration area (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"043", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"008", x"033", x"100");
	-- Test Case 19.6 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 0 Bytes from AEB3 critical configuration area (0x00040014)
	constant c_RMAP_CMD_TEST_CASE_19_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"044", x"000", x"000", x"004", x"000", x"014", x"000", x"000", x"000", x"0F9", x"100");
	-- Test Case 19.7 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"045", x"000", x"000", x"004", x"001", x"030", x"000", x"000", x"004", x"028", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 19.8 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 256 Bytes to AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_08_DATA : t_rmap_cmd_274_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"046", x"000", x"000", x"004", x"001", x"030", x"000", x"001", x"000", x"036", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"0A9", x"100");
	-- Test Case 19.9 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 260 Bytes to AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_09_DATA : t_rmap_cmd_278_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"047", x"000", x"000", x"004", x"001", x"030", x"000", x"001", x"004", x"01D", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"018", x"100");
	-- Test Case 19.10 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_10_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"048", x"000", x"000", x"004", x"001", x"030", x"000", x"000", x"000", x"012", x"000", x"100");
	-- Test Case 19.11 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"049", x"000", x"000", x"004", x"001", x"030", x"000", x"000", x"004", x"043", x"100");
	-- Test Case 19.12 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04A", x"000", x"000", x"004", x"001", x"030", x"000", x"001", x"000", x"05D", x"100");
	-- Test Case 19.13 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_13_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04B", x"000", x"000", x"004", x"001", x"030", x"000", x"001", x"004", x"076", x"100");
	-- Test Case 19.14 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB3 general configuration area (0x00040130)
	constant c_RMAP_CMD_TEST_CASE_19_14_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04C", x"000", x"000", x"004", x"001", x"030", x"000", x"000", x"000", x"0D8", x"100");
	-- Test Case 19.15 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB3 housekeeping area (0x00041000)
	constant c_RMAP_CMD_TEST_CASE_19_15_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04D", x"000", x"000", x"004", x"010", x"000", x"000", x"000", x"004", x"095", x"100");
	-- Test Case 19.16 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB3 housekeeping area (0x00041000)
	constant c_RMAP_CMD_TEST_CASE_19_16_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04E", x"000", x"000", x"004", x"010", x"000", x"000", x"001", x"000", x"08B", x"100");
	-- Test Case 19.17 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB3 housekeeping area (0x00041000)
	constant c_RMAP_CMD_TEST_CASE_19_17_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"04F", x"000", x"000", x"004", x"010", x"000", x"000", x"001", x"004", x"0A0", x"100");
	-- Test Case 19.18 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB3 housekeeping area (0x00041000)
	constant c_RMAP_CMD_TEST_CASE_19_18_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"050", x"000", x"000", x"004", x"010", x"000", x"000", x"000", x"000", x"02C", x"100");
	-- Test Case 20.1 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 bytes to AEB4 critical configuration are (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_01_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"051", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"004", x"003", x"000", x"000", x"000", x"0EE", x"042", x"100");
	-- Test Case 20.2 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 8 Bytes to AEB4 critical configuration area (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_02_DATA : t_rmap_cmd_26_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"052", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"008", x"07E", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"0FF", x"100");
	-- Test Case 20.3 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB4 critical configuration area (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_03_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"07C", x"0D1", x"050", x"000", x"053", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"000", x"05C", x"000", x"100");
	-- Test Case 20.4 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 4 Bytes from AEB4 critical configuration area (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_04_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"054", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"004", x"0D8", x"100");
	-- Test Case 20.5 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 8 Bytes from AEB4 critical configuration area (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_05_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"055", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"008", x"0FD", x"100");
	-- Test Case 20.6 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Read 0 Bytes from AEB4 critical configuration area (0x00080014)
	constant c_RMAP_CMD_TEST_CASE_20_06_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"056", x"000", x"000", x"008", x"000", x"014", x"000", x"000", x"000", x"087", x"100");
	-- Test Case 20.7 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 4 Bytes to AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_07_DATA : t_rmap_cmd_22_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"057", x"000", x"000", x"008", x"001", x"030", x"000", x"000", x"004", x"056", x"011", x"022", x"033", x"044", x"0CA", x"100");
	-- Test Case 20.8 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 256 Bytes to AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_08_DATA : t_rmap_cmd_274_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"058", x"000", x"000", x"008", x"001", x"030", x"000", x"001", x"000", x"059", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"0A9", x"100");
	-- Test Case 20.9 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 260 Bytes to AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_09_DATA : t_rmap_cmd_278_data  := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"059", x"000", x"000", x"008", x"001", x"030", x"000", x"001", x"004", x"072", x"011", x"022", x"033", x"044", x"055", x"066", x"077", x"088", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"018", x"100");
	-- Test Case 20.10 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Writing 0 Bytes to AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_10_DATA : t_rmap_cmd_18_data   := (x"051", x"001", x"06C", x"0D1", x"050", x"000", x"05A", x"000", x"000", x"008", x"001", x"030", x"000", x"000", x"000", x"06C", x"000", x"100");
	-- Test Case 20.11 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_11_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"05B", x"000", x"000", x"008", x"001", x"030", x"000", x"000", x"004", x"03D", x"100");
	-- Test Case 20.12 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_12_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"05C", x"000", x"000", x"008", x"001", x"030", x"000", x"001", x"000", x"093", x"100");
	-- Test Case 20.13 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_13_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"05D", x"000", x"000", x"008", x"001", x"030", x"000", x"001", x"004", x"0B8", x"100");
	-- Test Case 20.14 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB4 general configuration area (0x00080130)
	constant c_RMAP_CMD_TEST_CASE_20_14_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"05E", x"000", x"000", x"008", x"001", x"030", x"000", x"000", x"000", x"0A6", x"100");
	-- Test Case 20.15 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 4 Bytes from AEB4 housekeeping area (0x00081000)
	constant c_RMAP_CMD_TEST_CASE_20_15_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"05F", x"000", x"000", x"008", x"010", x"000", x"000", x"000", x"004", x"0EB", x"100");
	-- Test Case 20.16 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 256 Bytes from AEB4 housekeeping area (0x00081000)
	constant c_RMAP_CMD_TEST_CASE_20_16_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"060", x"000", x"000", x"008", x"010", x"000", x"000", x"001", x"000", x"0A0", x"100");
	-- Test Case 20.17 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 260 Bytes from AEB4 housekeeping area (0x00081000)
	constant c_RMAP_CMD_TEST_CASE_20_17_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"061", x"000", x"000", x"008", x"010", x"000", x"000", x"001", x"004", x"08B", x"100");
	-- Test Case 20.18 (PLATO-DLR-PL-ICD-0007 4.5.1.12): Reading 0 Bytes from AEB4 housekeeping area (0x00081000)
	constant c_RMAP_CMD_TEST_CASE_20_18_DATA : t_rmap_cmd_17_data   := (x"051", x"001", x"04C", x"0D1", x"050", x"000", x"062", x"000", x"000", x"008", x"010", x"000", x"000", x"000", x"000", x"095", x"100");

end package rmap_tb_stimulli_cmd_pkg;

package body rmap_tb_stimulli_cmd_pkg is

end package body rmap_tb_stimulli_cmd_pkg;
