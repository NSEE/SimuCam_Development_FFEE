library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ftdi_protocol_pkg.all;

entity usb3_fifo_master_stimuli is
	port(
		clk_i                : in    std_logic;
		rst_i                : in    std_logic;
		umft_wr_n_pin_i      : in    std_logic                     := '1';
		umft_rd_n_pin_i      : in    std_logic                     := '1';
		umft_oe_n_pin_i      : in    std_logic                     := '1';
		umft_data_bus_io     : inout std_logic_vector(31 downto 0) := (others => 'Z');
		umft_wakeup_n_pin_io : inout std_logic                     := 'Z';
		umft_be_bus_io       : inout std_logic_vector(3 downto 0)  := (others => 'Z');
		umft_gpio_bus_io     : inout std_logic_vector(1 downto 0)  := (others => 'Z');
		umft_rxf_n_pin_o     : out   std_logic;
		umft_txe_n_pin_o     : out   std_logic
	);
end entity usb3_fifo_master_stimuli;

architecture RTL of usb3_fifo_master_stimuli is

	signal s_umft601a_data_out     : std_logic_vector(31 downto 0);
	signal s_umft601a_wakeup_n_out : std_logic;
	signal s_umft601a_be_out       : std_logic_vector(3 downto 0);
	signal s_umft601a_gpio_out     : std_logic_vector(1 downto 0);
	signal s_umft601a_oe           : std_logic;
	signal s_umft601a_data_in      : std_logic_vector(31 downto 0);
	signal s_umft601a_wakeup_n_in  : std_logic;
	signal s_umft601a_be_in        : std_logic_vector(3 downto 0);
	signal s_umft601a_gpio_in      : std_logic_vector(1 downto 0);

	signal s_counter   : natural := 0;
	signal s_counter2  : natural := 0;
	signal s_times_cnt : natural := 0;

	-- ACK Package
	type t_ftdi_prot_ack_package is array (0 to 7) of std_logic_vector(31 downto 0);
	constant c_FTDI_PROT_ACK_PACKAGE  : t_ftdi_prot_ack_package := (
		c_FTDI_PROT_START_OF_PACKAGE,
		c_FTDI_PROT_PKG_ID_ACK_OK,
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"58374840",
		c_FTDI_PROT_END_OF_HEADER
	);
	constant c_FTDI_PROT_NACK_PACKAGE : t_ftdi_prot_ack_package := (
		c_FTDI_PROT_START_OF_PACKAGE,
		c_FTDI_PROT_PKG_ID_NACK_ERROR,
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"C7CEA3C5",
		c_FTDI_PROT_END_OF_HEADER
	);

	-- Reply Package
	type t_ftdi_prot_reply_package is array (0 to 7) of std_logic_vector(31 downto 0);
	constant c_FTDI_PROT_REPLY_PACKAGE : t_ftdi_prot_reply_package := (
		c_FTDI_PROT_START_OF_PACKAGE,
		c_FTDI_PROT_PKG_ID_HALF_CCD_REPLY,
		x"01020300",
		x"07001000",
		x"6B030000",
		x"008A0000",
		x"D48A4F2E",
		c_FTDI_PROT_END_OF_HEADER
	);

	-- Reply Payload
	type t_ftdi_prot_reply_payload is array (0 to 8834) of std_logic_vector(31 downto 0);
	constant c_FTDI_PROT_REPLY_PAYLOAD : t_ftdi_prot_reply_payload := (
		c_FTDI_PROT_START_OF_PAYLOAD,
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"00000100", x"02000300", x"04000500", x"06000700", x"08000900", x"0A000B00", x"0C000D00", x"0E000F00",
		x"10001100", x"12001300", x"14001500", x"16001700", x"18001900", x"1A001B00", x"1C001D00", x"1E001F00",
		x"20002100", x"22002300", x"24002500", x"26002700", x"28002900", x"2A002B00", x"2C002D00", x"2E002F00",
		x"30003100", x"32003300", x"34003500", x"36003700", x"38003900", x"3A003B00", x"3C003D00", x"3E003F00",
		x"FFFFFFFF", x"FFFFFFFF", x"40004100", x"42004300", x"44004500", x"46004700", x"48004900", x"4A004B00",
		x"4C004D00", x"4E004F00", x"50005100", x"52005300", x"54005500", x"56005700", x"58005900", x"5A005B00",
		x"5C005D00", x"5E005F00", x"60006100", x"62006300", x"64006500", x"66006700", x"68006900", x"6A006B00",
		x"6C006D00", x"6E006F00", x"70007100", x"72007300", x"74007500", x"76007700", x"78007900", x"7A007B00",
		x"7C007D00", x"7E007F00", x"FFFFFFFF", x"FFFFFFFF", x"80008100", x"82008300", x"84008500", x"86008700",
		x"88008900", x"8A008B00", x"8C008D00", x"8E008F00", x"90009100", x"92009300", x"94009500", x"96009700",
		x"98009900", x"9A009B00", x"9C009D00", x"9E009F00", x"A000A100", x"A200A300", x"A400A500", x"A600A700",
		x"A800A900", x"AA00AB00", x"AC00AD00", x"AE00AF00", x"B000B100", x"B200B300", x"B400B500", x"B600B700",
		x"B800B900", x"BA00BB00", x"BC00BD00", x"BE00BF00", x"FFFFFFFF", x"FFFFFFFF", x"C000C100", x"C200C300",
		x"C400C500", x"C600C700", x"C800C900", x"CA00CB00", x"CC00CD00", x"CE00CF00", x"D000D100", x"D200D300",
		x"D400D500", x"D600D700", x"D800D900", x"DA00DB00", x"DC00DD00", x"DE00DF00", x"E000E100", x"E200E300",
		x"E400E500", x"E600E700", x"E800E900", x"EA00EB00", x"EC00ED00", x"EE00EF00", x"F000F100", x"F200F300",
		x"F400F500", x"F600F700", x"F800F900", x"FA00FB00", x"FC00FD00", x"FE00FF00", x"FFFFFFFF", x"FFFFFFFF",
		x"00010101", x"02010301", x"04010501", x"06010701", x"08010901", x"0A010B01", x"0C010D01", x"0E010F01",
		x"10011101", x"12011301", x"14011501", x"16011701", x"18011901", x"1A011B01", x"1C011D01", x"1E011F01",
		x"20012101", x"22012301", x"24012501", x"26012701", x"28012901", x"2A012B01", x"2C012D01", x"2E012F01",
		x"30013101", x"32013301", x"34013501", x"36013701", x"38013901", x"3A013B01", x"3C013D01", x"3E013F01",
		x"FFFFFFFF", x"FFFFFFFF", x"40014101", x"42014301", x"44014501", x"46014701", x"48014901", x"4A014B01",
		x"4C014D01", x"4E014F01", x"50015101", x"52015301", x"54015501", x"56015701", x"58015901", x"5A015B01",
		x"5C015D01", x"5E015F01", x"60016101", x"62016301", x"64016501", x"66016701", x"68016901", x"6A016B01",
		x"6C016D01", x"6E016F01", x"70017101", x"72017301", x"74017501", x"76017701", x"78017901", x"7A017B01",
		x"7C017D01", x"7E017F01", x"FFFFFFFF", x"FFFFFFFF", x"80018101", x"82018301", x"84018501", x"86018701",
		x"88018901", x"8A018B01", x"8C018D01", x"8E018F01", x"90019101", x"92019301", x"94019501", x"96019701",
		x"98019901", x"9A019B01", x"9C019D01", x"9E019F01", x"A001A101", x"A201A301", x"A401A501", x"A601A701",
		x"A801A901", x"AA01AB01", x"AC01AD01", x"AE01AF01", x"B001B101", x"B201B301", x"B401B501", x"B601B701",
		x"B801B901", x"BA01BB01", x"BC01BD01", x"BE01BF01", x"FFFFFFFF", x"FFFFFFFF", x"C001C101", x"C201C301",
		x"C401C501", x"C601C701", x"C801C901", x"CA01CB01", x"CC01CD01", x"CE01CF01", x"D001D101", x"D201D301",
		x"D401D501", x"D601D701", x"D801D901", x"DA01DB01", x"DC01DD01", x"DE01DF01", x"E001E101", x"E201E301",
		x"E401E501", x"E601E701", x"E801E901", x"EA01EB01", x"EC01ED01", x"EE01EF01", x"F001F101", x"F201F301",
		x"F401F501", x"F601F701", x"F801F901", x"FA01FB01", x"FC01FD01", x"FE01FF01", x"FFFFFFFF", x"FFFFFFFF",
		x"00020102", x"02020302", x"04020502", x"06020702", x"08020902", x"0A020B02", x"0C020D02", x"0E020F02",
		x"10021102", x"12021302", x"14021502", x"16021702", x"18021902", x"1A021B02", x"1C021D02", x"1E021F02",
		x"20022102", x"22022302", x"24022502", x"26022702", x"28022902", x"2A022B02", x"2C022D02", x"2E022F02",
		x"30023102", x"32023302", x"34023502", x"36023702", x"38023902", x"3A023B02", x"3C023D02", x"3E023F02",
		x"FFFFFFFF", x"FFFFFFFF", x"40024102", x"42024302", x"44024502", x"46024702", x"48024902", x"4A024B02",
		x"4C024D02", x"4E024F02", x"50025102", x"52025302", x"54025502", x"56025702", x"58025902", x"5A025B02",
		x"5C025D02", x"5E025F02", x"60026102", x"62026302", x"64026502", x"66026702", x"68026902", x"6A026B02",
		x"6C026D02", x"6E026F02", x"70027102", x"72027302", x"74027502", x"76027702", x"78027902", x"7A027B02",
		x"7C027D02", x"7E027F02", x"FFFFFFFF", x"FFFFFFFF", x"80028102", x"82028302", x"84028502", x"86028702",
		x"88028902", x"8A028B02", x"8C028D02", x"8E028F02", x"90029102", x"92029302", x"94029502", x"96029702",
		x"98029902", x"9A029B02", x"9C029D02", x"9E029F02", x"A002A102", x"A202A302", x"A402A502", x"A602A702",
		x"A802A902", x"AA02AB02", x"AC02AD02", x"AE02AF02", x"B002B102", x"B202B302", x"B402B502", x"B602B702",
		x"B802B902", x"BA02BB02", x"BC02BD02", x"BE02BF02", x"FFFFFFFF", x"FFFFFFFF", x"C002C102", x"C202C302",
		x"C402C502", x"C602C702", x"C802C902", x"CA02CB02", x"CC02CD02", x"CE02CF02", x"D002D102", x"D202D302",
		x"D402D502", x"D602D702", x"D802D902", x"DA02DB02", x"DC02DD02", x"DE02DF02", x"E002E102", x"E202E302",
		x"E402E502", x"E602E702", x"E802E902", x"EA02EB02", x"EC02ED02", x"EE02EF02", x"F002F102", x"F202F302",
		x"F402F502", x"F602F702", x"F802F902", x"FA02FB02", x"FC02FD02", x"FE02FF02", x"FFFFFFFF", x"FFFFFFFF",
		x"00030103", x"02030303", x"04030503", x"06030703", x"08030903", x"0A030B03", x"0C030D03", x"0E030F03",
		x"10031103", x"12031303", x"14031503", x"16031703", x"18031903", x"1A031B03", x"1C031D03", x"1E031F03",
		x"20032103", x"22032303", x"24032503", x"26032703", x"28032903", x"2A032B03", x"2C032D03", x"2E032F03",
		x"30033103", x"32033303", x"34033503", x"36033703", x"38033903", x"3A033B03", x"3C033D03", x"3E033F03",
		x"FFFFFFFF", x"FFFFFFFF", x"40034103", x"42034303", x"44034503", x"46034703", x"48034903", x"4A034B03",
		x"4C034D03", x"4E034F03", x"50035103", x"52035303", x"54035503", x"56035703", x"58035903", x"5A035B03",
		x"5C035D03", x"5E035F03", x"60036103", x"62036303", x"64036503", x"66036703", x"68036903", x"6A036B03",
		x"6C036D03", x"6E036F03", x"70037103", x"72037303", x"74037503", x"76037703", x"78037903", x"7A037B03",
		x"7C037D03", x"7E037F03", x"FFFFFFFF", x"FFFFFFFF", x"80038103", x"82038303", x"84038503", x"86038703",
		x"88038903", x"8A038B03", x"8C038D03", x"8E038F03", x"90039103", x"92039303", x"94039503", x"96039703",
		x"98039903", x"9A039B03", x"9C039D03", x"9E039F03", x"A003A103", x"A203A303", x"A403A503", x"A603A703",
		x"A803A903", x"AA03AB03", x"AC03AD03", x"AE03AF03", x"B003B103", x"B203B303", x"B403B503", x"B603B703",
		x"B803B903", x"BA03BB03", x"BC03BD03", x"BE03BF03", x"FFFFFFFF", x"FFFFFFFF", x"C003C103", x"C203C303",
		x"C403C503", x"C603C703", x"C803C903", x"CA03CB03", x"CC03CD03", x"CE03CF03", x"D003D103", x"D203D303",
		x"D403D503", x"D603D703", x"D803D903", x"DA03DB03", x"DC03DD03", x"DE03DF03", x"E003E103", x"E203E303",
		x"E403E503", x"E603E703", x"E803E903", x"EA03EB03", x"EC03ED03", x"EE03EF03", x"F003F103", x"F203F303",
		x"F403F503", x"F603F703", x"F803F903", x"FA03FB03", x"FC03FD03", x"FE03FF03", x"FFFFFFFF", x"FFFFFFFF",
		x"00040104", x"02040304", x"04040504", x"06040704", x"08040904", x"0A040B04", x"0C040D04", x"0E040F04",
		x"10041104", x"12041304", x"14041504", x"16041704", x"18041904", x"1A041B04", x"1C041D04", x"1E041F04",
		x"20042104", x"22042304", x"24042504", x"26042704", x"28042904", x"2A042B04", x"2C042D04", x"2E042F04",
		x"30043104", x"32043304", x"34043504", x"36043704", x"38043904", x"3A043B04", x"3C043D04", x"3E043F04",
		x"FFFFFFFF", x"FFFFFFFF", x"40044104", x"42044304", x"44044504", x"46044704", x"48044904", x"4A044B04",
		x"4C044D04", x"4E044F04", x"50045104", x"52045304", x"54045504", x"56045704", x"58045904", x"5A045B04",
		x"5C045D04", x"5E045F04", x"60046104", x"62046304", x"64046504", x"66046704", x"68046904", x"6A046B04",
		x"6C046D04", x"6E046F04", x"70047104", x"72047304", x"74047504", x"76047704", x"78047904", x"7A047B04",
		x"7C047D04", x"7E047F04", x"FFFFFFFF", x"FFFFFFFF", x"80048104", x"82048304", x"84048504", x"86048704",
		x"88048904", x"8A048B04", x"8C048D04", x"8E048F04", x"90049104", x"92049304", x"94049504", x"96049704",
		x"98049904", x"9A049B04", x"9C049D04", x"9E049F04", x"A004A104", x"A204A304", x"A404A504", x"A604A704",
		x"A804A904", x"AA04AB04", x"AC04AD04", x"AE04AF04", x"B004B104", x"B204B304", x"B404B504", x"B604B704",
		x"B804B904", x"BA04BB04", x"BC04BD04", x"BE04BF04", x"FFFFFFFF", x"FFFFFFFF", x"C004C104", x"C204C304",
		x"C404C504", x"C604C704", x"C804C904", x"CA04CB04", x"CC04CD04", x"CE04CF04", x"D004D104", x"D204D304",
		x"D404D504", x"D604D704", x"D804D904", x"DA04DB04", x"DC04DD04", x"DE04DF04", x"E004E104", x"E204E304",
		x"E404E504", x"E604E704", x"E804E904", x"EA04EB04", x"EC04ED04", x"EE04EF04", x"F004F104", x"F204F304",
		x"F404F504", x"F604F704", x"F804F904", x"FA04FB04", x"FC04FD04", x"FE04FF04", x"FFFFFFFF", x"FFFFFFFF",
		x"00050105", x"02050305", x"04050505", x"06050705", x"08050905", x"0A050B05", x"0C050D05", x"0E050F05",
		x"10051105", x"12051305", x"14051505", x"16051705", x"18051905", x"1A051B05", x"1C051D05", x"1E051F05",
		x"20052105", x"22052305", x"24052505", x"26052705", x"28052905", x"2A052B05", x"2C052D05", x"2E052F05",
		x"30053105", x"32053305", x"34053505", x"36053705", x"38053905", x"3A053B05", x"3C053D05", x"3E053F05",
		x"FFFFFFFF", x"FFFFFFFF", x"40054105", x"42054305", x"44054505", x"46054705", x"48054905", x"4A054B05",
		x"4C054D05", x"4E054F05", x"50055105", x"52055305", x"54055505", x"56055705", x"58055905", x"5A055B05",
		x"5C055D05", x"5E055F05", x"60056105", x"62056305", x"64056505", x"66056705", x"68056905", x"6A056B05",
		x"6C056D05", x"6E056F05", x"70057105", x"72057305", x"74057505", x"76057705", x"78057905", x"7A057B05",
		x"7C057D05", x"7E057F05", x"FFFFFFFF", x"FFFFFFFF", x"80058105", x"82058305", x"84058505", x"86058705",
		x"88058905", x"8A058B05", x"8C058D05", x"8E058F05", x"90059105", x"92059305", x"94059505", x"96059705",
		x"98059905", x"9A059B05", x"9C059D05", x"9E059F05", x"A005A105", x"A205A305", x"A405A505", x"A605A705",
		x"A805A905", x"AA05AB05", x"AC05AD05", x"AE05AF05", x"B005B105", x"B205B305", x"B405B505", x"B605B705",
		x"B805B905", x"BA05BB05", x"BC05BD05", x"BE05BF05", x"FFFFFFFF", x"FFFFFFFF", x"C005C105", x"C205C305",
		x"C405C505", x"C605C705", x"C805C905", x"CA05CB05", x"CC05CD05", x"CE05CF05", x"D005D105", x"D205D305",
		x"D405D505", x"D605D705", x"D805D905", x"DA05DB05", x"DC05DD05", x"DE05DF05", x"E005E105", x"E205E305",
		x"E405E505", x"E605E705", x"E805E905", x"EA05EB05", x"EC05ED05", x"EE05EF05", x"F005F105", x"F205F305",
		x"F405F505", x"F605F705", x"F805F905", x"FA05FB05", x"FC05FD05", x"FE05FF05", x"FFFFFFFF", x"FFFFFFFF",
		x"00060106", x"02060306", x"04060506", x"06060706", x"08060906", x"0A060B06", x"0C060D06", x"0E060F06",
		x"10061106", x"12061306", x"14061506", x"16061706", x"18061906", x"1A061B06", x"1C061D06", x"1E061F06",
		x"20062106", x"22062306", x"24062506", x"26062706", x"28062906", x"2A062B06", x"2C062D06", x"2E062F06",
		x"30063106", x"32063306", x"34063506", x"36063706", x"38063906", x"3A063B06", x"3C063D06", x"3E063F06",
		x"FFFFFFFF", x"FFFFFFFF", x"40064106", x"42064306", x"44064506", x"46064706", x"48064906", x"4A064B06",
		x"4C064D06", x"4E064F06", x"50065106", x"52065306", x"54065506", x"56065706", x"58065906", x"5A065B06",
		x"5C065D06", x"5E065F06", x"60066106", x"62066306", x"64066506", x"66066706", x"68066906", x"6A066B06",
		x"6C066D06", x"6E066F06", x"70067106", x"72067306", x"74067506", x"76067706", x"78067906", x"7A067B06",
		x"7C067D06", x"7E067F06", x"FFFFFFFF", x"FFFFFFFF", x"80068106", x"82068306", x"84068506", x"86068706",
		x"88068906", x"8A068B06", x"8C068D06", x"8E068F06", x"90069106", x"92069306", x"94069506", x"96069706",
		x"98069906", x"9A069B06", x"9C069D06", x"9E069F06", x"A006A106", x"A206A306", x"A406A506", x"A606A706",
		x"A806A906", x"AA06AB06", x"AC06AD06", x"AE06AF06", x"B006B106", x"B206B306", x"B406B506", x"B606B706",
		x"B806B906", x"BA06BB06", x"BC06BD06", x"BE06BF06", x"FFFFFFFF", x"FFFFFFFF", x"C006C106", x"C206C306",
		x"C406C506", x"C606C706", x"C806C906", x"CA06CB06", x"CC06CD06", x"CE06CF06", x"D006D106", x"D206D306",
		x"D406D506", x"D606D706", x"D806D906", x"DA06DB06", x"DC06DD06", x"DE06DF06", x"E006E106", x"E206E306",
		x"E406E506", x"E606E706", x"E806E906", x"EA06EB06", x"EC06ED06", x"EE06EF06", x"F006F106", x"F206F306",
		x"F406F506", x"F606F706", x"F806F906", x"FA06FB06", x"FC06FD06", x"FE06FF06", x"FFFFFFFF", x"FFFFFFFF",
		x"00070107", x"02070307", x"04070507", x"06070707", x"08070907", x"0A070B07", x"0C070D07", x"0E070F07",
		x"10071107", x"12071307", x"14071507", x"16071707", x"18071907", x"1A071B07", x"1C071D07", x"1E071F07",
		x"20072107", x"22072307", x"24072507", x"26072707", x"28072907", x"2A072B07", x"2C072D07", x"2E072F07",
		x"30073107", x"32073307", x"34073507", x"36073707", x"38073907", x"3A073B07", x"3C073D07", x"3E073F07",
		x"FFFFFFFF", x"FFFFFFFF", x"40074107", x"42074307", x"44074507", x"46074707", x"48074907", x"4A074B07",
		x"4C074D07", x"4E074F07", x"50075107", x"52075307", x"54075507", x"56075707", x"58075907", x"5A075B07",
		x"5C075D07", x"5E075F07", x"60076107", x"62076307", x"64076507", x"66076707", x"68076907", x"6A076B07",
		x"6C076D07", x"6E076F07", x"70077107", x"72077307", x"74077507", x"76077707", x"78077907", x"7A077B07",
		x"7C077D07", x"7E077F07", x"FFFFFFFF", x"FFFFFFFF", x"80078107", x"82078307", x"84078507", x"86078707",
		x"88078907", x"8A078B07", x"8C078D07", x"8E078F07", x"90079107", x"92079307", x"94079507", x"96079707",
		x"98079907", x"9A079B07", x"9C079D07", x"9E079F07", x"A007A107", x"A207A307", x"A407A507", x"A607A707",
		x"A807A907", x"AA07AB07", x"AC07AD07", x"AE07AF07", x"B007B107", x"B207B307", x"B407B507", x"B607B707",
		x"B807B907", x"BA07BB07", x"BC07BD07", x"BE07BF07", x"FFFFFFFF", x"FFFFFFFF", x"C007C107", x"C207C307",
		x"C407C507", x"C607C707", x"C807C907", x"CA07CB07", x"CC07CD07", x"CE07CF07", x"D007D107", x"D207D307",
		x"D407D507", x"D607D707", x"D807D907", x"DA07DB07", x"DC07DD07", x"DE07DF07", x"E007E107", x"E207E307",
		x"E407E507", x"E607E707", x"E807E907", x"EA07EB07", x"EC07ED07", x"EE07EF07", x"F007F107", x"F207F307",
		x"F407F507", x"F607F707", x"F807F907", x"FA07FB07", x"FC07FD07", x"FE07FF07", x"FFFFFFFF", x"FFFFFFFF",
		x"00080108", x"02080308", x"04080508", x"06080708", x"08080908", x"0A080B08", x"0C080D08", x"0E080F08",
		x"10081108", x"12081308", x"14081508", x"16081708", x"18081908", x"1A081B08", x"1C081D08", x"1E081F08",
		x"20082108", x"22082308", x"24082508", x"26082708", x"28082908", x"2A082B08", x"2C082D08", x"2E082F08",
		x"30083108", x"32083308", x"34083508", x"36083708", x"38083908", x"3A083B08", x"3C083D08", x"3E083F08",
		x"FFFFFFFF", x"FFFFFFFF", x"40084108", x"42084308", x"44084508", x"46084708", x"48084908", x"4A084B08",
		x"4C084D08", x"4E084F08", x"50085108", x"52085308", x"54085508", x"56085708", x"58085908", x"5A085B08",
		x"5C085D08", x"5E085F08", x"60086108", x"62086308", x"64086508", x"66086708", x"68086908", x"6A086B08",
		x"6C086D08", x"6E086F08", x"70087108", x"72087308", x"74087508", x"76087708", x"78087908", x"7A087B08",
		x"7C087D08", x"7E087F08", x"FFFFFFFF", x"FFFFFFFF", x"80088108", x"82088308", x"84088508", x"86088708",
		x"88088908", x"8A088B08", x"8C088D08", x"8E088F08", x"90089108", x"92089308", x"94089508", x"96089708",
		x"98089908", x"9A089B08", x"9C089D08", x"9E089F08", x"A008A108", x"A208A308", x"A408A508", x"A608A708",
		x"A808A908", x"AA08AB08", x"AC08AD08", x"AE08AF08", x"B008B108", x"B208B308", x"B408B508", x"B608B708",
		x"B808B908", x"BA08BB08", x"BC08BD08", x"BE08BF08", x"FFFFFFFF", x"FFFFFFFF", x"C008C108", x"C208C308",
		x"C408C508", x"C608C708", x"C808C908", x"CA08CB08", x"CC08CD08", x"CE08CF08", x"D008D108", x"D208D308",
		x"D408D508", x"D608D708", x"D808D908", x"DA08DB08", x"DC08DD08", x"DE08DF08", x"E008E108", x"E208E308",
		x"E408E508", x"E608E708", x"E808E908", x"EA08EB08", x"EC08ED08", x"EE08EF08", x"F008F108", x"F208F308",
		x"F408F508", x"F608F708", x"F808F908", x"FA08FB08", x"FC08FD08", x"FE08FF08", x"FFFFFFFF", x"FFFFFFFF",
		x"00090109", x"02090309", x"04090509", x"06090709", x"08090909", x"0A090B09", x"0C090D09", x"0E090F09",
		x"10091109", x"12091309", x"14091509", x"16091709", x"18091909", x"1A091B09", x"1C091D09", x"1E091F09",
		x"20092109", x"22092309", x"24092509", x"26092709", x"28092909", x"2A092B09", x"2C092D09", x"2E092F09",
		x"30093109", x"32093309", x"34093509", x"36093709", x"38093909", x"3A093B09", x"3C093D09", x"3E093F09",
		x"FFFFFFFF", x"FFFFFFFF", x"40094109", x"42094309", x"44094509", x"46094709", x"48094909", x"4A094B09",
		x"4C094D09", x"4E094F09", x"50095109", x"52095309", x"54095509", x"56095709", x"58095909", x"5A095B09",
		x"5C095D09", x"5E095F09", x"60096109", x"62096309", x"64096509", x"66096709", x"68096909", x"6A096B09",
		x"6C096D09", x"6E096F09", x"70097109", x"72097309", x"74097509", x"76097709", x"78097909", x"7A097B09",
		x"7C097D09", x"7E097F09", x"FFFFFFFF", x"FFFFFFFF", x"80098109", x"82098309", x"84098509", x"86098709",
		x"88098909", x"8A098B09", x"8C098D09", x"8E098F09", x"90099109", x"92099309", x"94099509", x"96099709",
		x"98099909", x"9A099B09", x"9C099D09", x"9E099F09", x"A009A109", x"A209A309", x"A409A509", x"A609A709",
		x"A809A909", x"AA09AB09", x"AC09AD09", x"AE09AF09", x"B009B109", x"B209B309", x"B409B509", x"B609B709",
		x"B809B909", x"BA09BB09", x"BC09BD09", x"BE09BF09", x"FFFFFFFF", x"FFFFFFFF", x"C009C109", x"C209C309",
		x"C409C509", x"C609C709", x"C809C909", x"CA09CB09", x"CC09CD09", x"CE09CF09", x"D009D109", x"D209D309",
		x"D409D509", x"D609D709", x"D809D909", x"DA09DB09", x"DC09DD09", x"DE09DF09", x"E009E109", x"E209E309",
		x"E409E509", x"E609E709", x"E809E909", x"EA09EB09", x"EC09ED09", x"EE09EF09", x"F009F109", x"F209F309",
		x"F409F509", x"F609F709", x"F809F909", x"FA09FB09", x"FC09FD09", x"FE09FF09", x"FFFFFFFF", x"FFFFFFFF",
		x"000A010A", x"020A030A", x"040A050A", x"060A070A", x"080A090A", x"0A0A0B0A", x"0C0A0D0A", x"0E0A0F0A",
		x"100A110A", x"120A130A", x"140A150A", x"160A170A", x"180A190A", x"1A0A1B0A", x"1C0A1D0A", x"1E0A1F0A",
		x"200A210A", x"220A230A", x"240A250A", x"260A270A", x"280A290A", x"2A0A2B0A", x"2C0A2D0A", x"2E0A2F0A",
		x"300A310A", x"320A330A", x"340A350A", x"360A370A", x"380A390A", x"3A0A3B0A", x"3C0A3D0A", x"3E0A3F0A",
		x"FFFFFFFF", x"FFFFFFFF", x"400A410A", x"420A430A", x"440A450A", x"460A470A", x"480A490A", x"4A0A4B0A",
		x"4C0A4D0A", x"4E0A4F0A", x"500A510A", x"520A530A", x"540A550A", x"560A570A", x"580A590A", x"5A0A5B0A",
		x"5C0A5D0A", x"5E0A5F0A", x"600A610A", x"620A630A", x"640A650A", x"660A670A", x"680A690A", x"6A0A6B0A",
		x"6C0A6D0A", x"6E0A6F0A", x"700A710A", x"720A730A", x"740A750A", x"760A770A", x"780A790A", x"7A0A7B0A",
		x"7C0A7D0A", x"7E0A7F0A", x"FFFFFFFF", x"FFFFFFFF", x"800A810A", x"820A830A", x"840A850A", x"860A870A",
		x"880A890A", x"8A0A8B0A", x"8C0A8D0A", x"8E0A8F0A", x"900A910A", x"920A930A", x"940A950A", x"960A970A",
		x"980A990A", x"9A0A9B0A", x"9C0A9D0A", x"9E0A9F0A", x"A00AA10A", x"A20AA30A", x"A40AA50A", x"A60AA70A",
		x"A80AA90A", x"AA0AAB0A", x"AC0AAD0A", x"AE0AAF0A", x"B00AB10A", x"B20AB30A", x"B40AB50A", x"B60AB70A",
		x"B80AB90A", x"BA0ABB0A", x"BC0ABD0A", x"BE0ABF0A", x"FFFFFFFF", x"FFFFFFFF", x"C00AC10A", x"C20AC30A",
		x"C40AC50A", x"C60AC70A", x"C80AC90A", x"CA0ACB0A", x"CC0ACD0A", x"CE0ACF0A", x"D00AD10A", x"D20AD30A",
		x"D40AD50A", x"D60AD70A", x"D80AD90A", x"DA0ADB0A", x"DC0ADD0A", x"DE0ADF0A", x"E00AE10A", x"E20AE30A",
		x"E40AE50A", x"E60AE70A", x"E80AE90A", x"EA0AEB0A", x"EC0AED0A", x"EE0AEF0A", x"F00AF10A", x"F20AF30A",
		x"F40AF50A", x"F60AF70A", x"F80AF90A", x"FA0AFB0A", x"FC0AFD0A", x"FE0AFF0A", x"FFFFFFFF", x"FFFFFFFF",
		x"000B010B", x"020B030B", x"040B050B", x"060B070B", x"080B090B", x"0A0B0B0B", x"0C0B0D0B", x"0E0B0F0B",
		x"100B110B", x"120B130B", x"140B150B", x"160B170B", x"180B190B", x"1A0B1B0B", x"1C0B1D0B", x"1E0B1F0B",
		x"200B210B", x"220B230B", x"240B250B", x"260B270B", x"280B290B", x"2A0B2B0B", x"2C0B2D0B", x"2E0B2F0B",
		x"300B310B", x"320B330B", x"340B350B", x"360B370B", x"380B390B", x"3A0B3B0B", x"3C0B3D0B", x"3E0B3F0B",
		x"FFFFFFFF", x"FFFFFFFF", x"400B410B", x"420B430B", x"440B450B", x"460B470B", x"480B490B", x"4A0B4B0B",
		x"4C0B4D0B", x"4E0B4F0B", x"500B510B", x"520B530B", x"540B550B", x"560B570B", x"580B590B", x"5A0B5B0B",
		x"5C0B5D0B", x"5E0B5F0B", x"600B610B", x"620B630B", x"640B650B", x"660B670B", x"680B690B", x"6A0B6B0B",
		x"6C0B6D0B", x"6E0B6F0B", x"700B710B", x"720B730B", x"740B750B", x"760B770B", x"780B790B", x"7A0B7B0B",
		x"7C0B7D0B", x"7E0B7F0B", x"FFFFFFFF", x"FFFFFFFF", x"800B810B", x"820B830B", x"840B850B", x"860B870B",
		x"880B890B", x"8A0B8B0B", x"8C0B8D0B", x"8E0B8F0B", x"900B910B", x"920B930B", x"940B950B", x"960B970B",
		x"980B990B", x"9A0B9B0B", x"9C0B9D0B", x"9E0B9F0B", x"A00BA10B", x"A20BA30B", x"A40BA50B", x"A60BA70B",
		x"A80BA90B", x"AA0BAB0B", x"AC0BAD0B", x"AE0BAF0B", x"B00BB10B", x"B20BB30B", x"B40BB50B", x"B60BB70B",
		x"B80BB90B", x"BA0BBB0B", x"BC0BBD0B", x"BE0BBF0B", x"FFFFFFFF", x"FFFFFFFF", x"C00BC10B", x"C20BC30B",
		x"C40BC50B", x"C60BC70B", x"C80BC90B", x"CA0BCB0B", x"CC0BCD0B", x"CE0BCF0B", x"D00BD10B", x"D20BD30B",
		x"D40BD50B", x"D60BD70B", x"D80BD90B", x"DA0BDB0B", x"DC0BDD0B", x"DE0BDF0B", x"E00BE10B", x"E20BE30B",
		x"E40BE50B", x"E60BE70B", x"E80BE90B", x"EA0BEB0B", x"EC0BED0B", x"EE0BEF0B", x"F00BF10B", x"F20BF30B",
		x"F40BF50B", x"F60BF70B", x"F80BF90B", x"FA0BFB0B", x"FC0BFD0B", x"FE0BFF0B", x"FFFFFFFF", x"FFFFFFFF",
		x"000C010C", x"020C030C", x"040C050C", x"060C070C", x"080C090C", x"0A0C0B0C", x"0C0C0D0C", x"0E0C0F0C",
		x"100C110C", x"120C130C", x"140C150C", x"160C170C", x"180C190C", x"1A0C1B0C", x"1C0C1D0C", x"1E0C1F0C",
		x"200C210C", x"220C230C", x"240C250C", x"260C270C", x"280C290C", x"2A0C2B0C", x"2C0C2D0C", x"2E0C2F0C",
		x"300C310C", x"320C330C", x"340C350C", x"360C370C", x"380C390C", x"3A0C3B0C", x"3C0C3D0C", x"3E0C3F0C",
		x"FFFFFFFF", x"FFFFFFFF", x"400C410C", x"420C430C", x"440C450C", x"460C470C", x"480C490C", x"4A0C4B0C",
		x"4C0C4D0C", x"4E0C4F0C", x"500C510C", x"520C530C", x"540C550C", x"560C570C", x"580C590C", x"5A0C5B0C",
		x"5C0C5D0C", x"5E0C5F0C", x"600C610C", x"620C630C", x"640C650C", x"660C670C", x"680C690C", x"6A0C6B0C",
		x"6C0C6D0C", x"6E0C6F0C", x"700C710C", x"720C730C", x"740C750C", x"760C770C", x"780C790C", x"7A0C7B0C",
		x"7C0C7D0C", x"7E0C7F0C", x"FFFFFFFF", x"FFFFFFFF", x"800C810C", x"820C830C", x"840C850C", x"860C870C",
		x"880C890C", x"8A0C8B0C", x"8C0C8D0C", x"8E0C8F0C", x"900C910C", x"920C930C", x"940C950C", x"960C970C",
		x"980C990C", x"9A0C9B0C", x"9C0C9D0C", x"9E0C9F0C", x"A00CA10C", x"A20CA30C", x"A40CA50C", x"A60CA70C",
		x"A80CA90C", x"AA0CAB0C", x"AC0CAD0C", x"AE0CAF0C", x"B00CB10C", x"B20CB30C", x"B40CB50C", x"B60CB70C",
		x"B80CB90C", x"BA0CBB0C", x"BC0CBD0C", x"BE0CBF0C", x"FFFFFFFF", x"FFFFFFFF", x"C00CC10C", x"C20CC30C",
		x"C40CC50C", x"C60CC70C", x"C80CC90C", x"CA0CCB0C", x"CC0CCD0C", x"CE0CCF0C", x"D00CD10C", x"D20CD30C",
		x"D40CD50C", x"D60CD70C", x"D80CD90C", x"DA0CDB0C", x"DC0CDD0C", x"DE0CDF0C", x"E00CE10C", x"E20CE30C",
		x"E40CE50C", x"E60CE70C", x"E80CE90C", x"EA0CEB0C", x"EC0CED0C", x"EE0CEF0C", x"F00CF10C", x"F20CF30C",
		x"F40CF50C", x"F60CF70C", x"F80CF90C", x"FA0CFB0C", x"FC0CFD0C", x"FE0CFF0C", x"FFFFFFFF", x"FFFFFFFF",
		x"000D010D", x"020D030D", x"040D050D", x"060D070D", x"080D090D", x"0A0D0B0D", x"0C0D0D0D", x"0E0D0F0D",
		x"100D110D", x"120D130D", x"140D150D", x"160D170D", x"180D190D", x"1A0D1B0D", x"1C0D1D0D", x"1E0D1F0D",
		x"200D210D", x"220D230D", x"240D250D", x"260D270D", x"280D290D", x"2A0D2B0D", x"2C0D2D0D", x"2E0D2F0D",
		x"300D310D", x"320D330D", x"340D350D", x"360D370D", x"380D390D", x"3A0D3B0D", x"3C0D3D0D", x"3E0D3F0D",
		x"FFFFFFFF", x"FFFFFFFF", x"400D410D", x"420D430D", x"440D450D", x"460D470D", x"480D490D", x"4A0D4B0D",
		x"4C0D4D0D", x"4E0D4F0D", x"500D510D", x"520D530D", x"540D550D", x"560D570D", x"580D590D", x"5A0D5B0D",
		x"5C0D5D0D", x"5E0D5F0D", x"600D610D", x"620D630D", x"640D650D", x"660D670D", x"680D690D", x"6A0D6B0D",
		x"6C0D6D0D", x"6E0D6F0D", x"700D710D", x"720D730D", x"740D750D", x"760D770D", x"780D790D", x"7A0D7B0D",
		x"7C0D7D0D", x"7E0D7F0D", x"FFFFFFFF", x"FFFFFFFF", x"800D810D", x"820D830D", x"840D850D", x"860D870D",
		x"880D890D", x"8A0D8B0D", x"8C0D8D0D", x"8E0D8F0D", x"900D910D", x"920D930D", x"940D950D", x"960D970D",
		x"980D990D", x"9A0D9B0D", x"9C0D9D0D", x"9E0D9F0D", x"A00DA10D", x"A20DA30D", x"A40DA50D", x"A60DA70D",
		x"A80DA90D", x"AA0DAB0D", x"AC0DAD0D", x"AE0DAF0D", x"B00DB10D", x"B20DB30D", x"B40DB50D", x"B60DB70D",
		x"B80DB90D", x"BA0DBB0D", x"BC0DBD0D", x"BE0DBF0D", x"FFFFFFFF", x"FFFFFFFF", x"C00DC10D", x"C20DC30D",
		x"C40DC50D", x"C60DC70D", x"C80DC90D", x"CA0DCB0D", x"CC0DCD0D", x"CE0DCF0D", x"D00DD10D", x"D20DD30D",
		x"D40DD50D", x"D60DD70D", x"D80DD90D", x"DA0DDB0D", x"DC0DDD0D", x"DE0DDF0D", x"E00DE10D", x"E20DE30D",
		x"E40DE50D", x"E60DE70D", x"E80DE90D", x"EA0DEB0D", x"EC0DED0D", x"EE0DEF0D", x"F00DF10D", x"F20DF30D",
		x"F40DF50D", x"F60DF70D", x"F80DF90D", x"FA0DFB0D", x"FC0DFD0D", x"FE0DFF0D", x"FFFFFFFF", x"FFFFFFFF",
		x"000E010E", x"020E030E", x"040E050E", x"060E070E", x"080E090E", x"0A0E0B0E", x"0C0E0D0E", x"0E0E0F0E",
		x"100E110E", x"120E130E", x"140E150E", x"160E170E", x"180E190E", x"1A0E1B0E", x"1C0E1D0E", x"1E0E1F0E",
		x"200E210E", x"220E230E", x"240E250E", x"260E270E", x"280E290E", x"2A0E2B0E", x"2C0E2D0E", x"2E0E2F0E",
		x"300E310E", x"320E330E", x"340E350E", x"360E370E", x"380E390E", x"3A0E3B0E", x"3C0E3D0E", x"3E0E3F0E",
		x"FFFFFFFF", x"FFFFFFFF", x"400E410E", x"420E430E", x"440E450E", x"460E470E", x"480E490E", x"4A0E4B0E",
		x"4C0E4D0E", x"4E0E4F0E", x"500E510E", x"520E530E", x"540E550E", x"560E570E", x"580E590E", x"5A0E5B0E",
		x"5C0E5D0E", x"5E0E5F0E", x"600E610E", x"620E630E", x"640E650E", x"660E670E", x"680E690E", x"6A0E6B0E",
		x"6C0E6D0E", x"6E0E6F0E", x"700E710E", x"720E730E", x"740E750E", x"760E770E", x"780E790E", x"7A0E7B0E",
		x"7C0E7D0E", x"7E0E7F0E", x"FFFFFFFF", x"FFFFFFFF", x"800E810E", x"820E830E", x"840E850E", x"860E870E",
		x"880E890E", x"8A0E8B0E", x"8C0E8D0E", x"8E0E8F0E", x"900E910E", x"920E930E", x"940E950E", x"960E970E",
		x"980E990E", x"9A0E9B0E", x"9C0E9D0E", x"9E0E9F0E", x"A00EA10E", x"A20EA30E", x"A40EA50E", x"A60EA70E",
		x"A80EA90E", x"AA0EAB0E", x"AC0EAD0E", x"AE0EAF0E", x"B00EB10E", x"B20EB30E", x"B40EB50E", x"B60EB70E",
		x"B80EB90E", x"BA0EBB0E", x"BC0EBD0E", x"BE0EBF0E", x"FFFFFFFF", x"FFFFFFFF", x"C00EC10E", x"C20EC30E",
		x"C40EC50E", x"C60EC70E", x"C80EC90E", x"CA0ECB0E", x"CC0ECD0E", x"CE0ECF0E", x"D00ED10E", x"D20ED30E",
		x"D40ED50E", x"D60ED70E", x"D80ED90E", x"DA0EDB0E", x"DC0EDD0E", x"DE0EDF0E", x"E00EE10E", x"E20EE30E",
		x"E40EE50E", x"E60EE70E", x"E80EE90E", x"EA0EEB0E", x"EC0EED0E", x"EE0EEF0E", x"F00EF10E", x"F20EF30E",
		x"F40EF50E", x"F60EF70E", x"F80EF90E", x"FA0EFB0E", x"FC0EFD0E", x"FE0EFF0E", x"FFFFFFFF", x"FFFFFFFF",
		x"000F010F", x"020F030F", x"040F050F", x"060F070F", x"080F090F", x"0A0F0B0F", x"0C0F0D0F", x"0E0F0F0F",
		x"100F110F", x"120F130F", x"140F150F", x"160F170F", x"180F190F", x"1A0F1B0F", x"1C0F1D0F", x"1E0F1F0F",
		x"200F210F", x"220F230F", x"240F250F", x"260F270F", x"280F290F", x"2A0F2B0F", x"2C0F2D0F", x"2E0F2F0F",
		x"300F310F", x"320F330F", x"340F350F", x"360F370F", x"380F390F", x"3A0F3B0F", x"3C0F3D0F", x"3E0F3F0F",
		x"FFFFFFFF", x"FFFFFFFF", x"400F410F", x"420F430F", x"440F450F", x"460F470F", x"480F490F", x"4A0F4B0F",
		x"4C0F4D0F", x"4E0F4F0F", x"500F510F", x"520F530F", x"540F550F", x"560F570F", x"580F590F", x"5A0F5B0F",
		x"5C0F5D0F", x"5E0F5F0F", x"600F610F", x"620F630F", x"640F650F", x"660F670F", x"680F690F", x"6A0F6B0F",
		x"6C0F6D0F", x"6E0F6F0F", x"700F710F", x"720F730F", x"740F750F", x"760F770F", x"780F790F", x"7A0F7B0F",
		x"7C0F7D0F", x"7E0F7F0F", x"FFFFFFFF", x"FFFFFFFF", x"800F810F", x"820F830F", x"840F850F", x"860F870F",
		x"880F890F", x"8A0F8B0F", x"8C0F8D0F", x"8E0F8F0F", x"900F910F", x"920F930F", x"940F950F", x"960F970F",
		x"980F990F", x"9A0F9B0F", x"9C0F9D0F", x"9E0F9F0F", x"A00FA10F", x"A20FA30F", x"A40FA50F", x"A60FA70F",
		x"A80FA90F", x"AA0FAB0F", x"AC0FAD0F", x"AE0FAF0F", x"B00FB10F", x"B20FB30F", x"B40FB50F", x"B60FB70F",
		x"B80FB90F", x"BA0FBB0F", x"BC0FBD0F", x"BE0FBF0F", x"FFFFFFFF", x"FFFFFFFF", x"C00FC10F", x"C20FC30F",
		x"C40FC50F", x"C60FC70F", x"C80FC90F", x"CA0FCB0F", x"CC0FCD0F", x"CE0FCF0F", x"D00FD10F", x"D20FD30F",
		x"D40FD50F", x"D60FD70F", x"D80FD90F", x"DA0FDB0F", x"DC0FDD0F", x"DE0FDF0F", x"E00FE10F", x"E20FE30F",
		x"E40FE50F", x"E60FE70F", x"E80FE90F", x"EA0FEB0F", x"EC0FED0F", x"EE0FEF0F", x"F00FF10F", x"F20FF30F",
		x"F40FF50F", x"F60FF70F", x"F80FF90F", x"FA0FFB0F", x"FC0FFD0F", x"FE0FFF0F", x"FFFFFFFF", x"FFFFFFFF",
		x"00100110", x"02100310", x"04100510", x"06100710", x"08100910", x"0A100B10", x"0C100D10", x"0E100F10",
		x"10101110", x"12101310", x"14101510", x"16101710", x"18101910", x"1A101B10", x"1C101D10", x"1E101F10",
		x"20102110", x"22102310", x"24102510", x"26102710", x"28102910", x"2A102B10", x"2C102D10", x"2E102F10",
		x"30103110", x"32103310", x"34103510", x"36103710", x"38103910", x"3A103B10", x"3C103D10", x"3E103F10",
		x"FFFFFFFF", x"FFFFFFFF", x"40104110", x"42104310", x"44104510", x"46104710", x"48104910", x"4A104B10",
		x"4C104D10", x"4E104F10", x"50105110", x"52105310", x"54105510", x"56105710", x"58105910", x"5A105B10",
		x"5C105D10", x"5E105F10", x"60106110", x"62106310", x"64106510", x"66106710", x"68106910", x"6A106B10",
		x"6C106D10", x"6E106F10", x"70107110", x"72107310", x"74107510", x"76107710", x"78107910", x"7A107B10",
		x"7C107D10", x"7E107F10", x"FFFFFFFF", x"FFFFFFFF", x"80108110", x"82108310", x"84108510", x"86108710",
		x"88108910", x"8A108B10", x"8C108D10", x"8E108F10", x"90109110", x"92109310", x"94109510", x"96109710",
		x"98109910", x"9A109B10", x"9C109D10", x"9E109F10", x"A010A110", x"A210A310", x"A410A510", x"A610A710",
		x"A810A910", x"AA10AB10", x"AC10AD10", x"AE10AF10", x"B010B110", x"B210B310", x"B410B510", x"B610B710",
		x"B810B910", x"BA10BB10", x"BC10BD10", x"BE10BF10", x"FFFFFFFF", x"FFFFFFFF", x"C010C110", x"C210C310",
		x"C410C510", x"C610C710", x"C810C910", x"CA10CB10", x"CC10CD10", x"CE10CF10", x"D010D110", x"D210D310",
		x"D410D510", x"D610D710", x"D810D910", x"DA10DB10", x"DC10DD10", x"DE10DF10", x"E010E110", x"E210E310",
		x"E410E510", x"E610E710", x"E810E910", x"EA10EB10", x"EC10ED10", x"EE10EF10", x"F010F110", x"F210F310",
		x"F410F510", x"F610F710", x"F810F910", x"FA10FB10", x"FC10FD10", x"FE10FF10", x"FFFFFFFF", x"FFFFFFFF",
		x"00110111", x"02110311", x"04110511", x"06110711", x"08110911", x"0A110B11", x"0C110D11", x"0E110F11",
		x"10111111", x"12111311", x"14111511", x"16111711", x"18111911", x"1A111B11", x"1C111D11", x"1E111F11",
		x"20112111", x"22112311", x"24112511", x"26112711", x"28112911", x"2A112B11", x"2C112D11", x"2E112F11",
		x"30113111", x"32113311", x"34113511", x"36113711", x"38113911", x"3A113B11", x"3C113D11", x"3E113F11",
		x"FFFFFFFF", x"FFFFFFFF", x"40114111", x"42114311", x"44114511", x"46114711", x"48114911", x"4A114B11",
		x"4C114D11", x"4E114F11", x"50115111", x"52115311", x"54115511", x"56115711", x"58115911", x"5A115B11",
		x"5C115D11", x"5E115F11", x"60116111", x"62116311", x"64116511", x"66116711", x"68116911", x"6A116B11",
		x"6C116D11", x"6E116F11", x"70117111", x"72117311", x"74117511", x"76117711", x"78117911", x"7A117B11",
		x"7C117D11", x"7E117F11", x"FFFFFFFF", x"FFFFFFFF", x"80118111", x"82118311", x"84118511", x"86118711",
		x"88118911", x"8A118B11", x"8C118D11", x"8E118F11", x"90119111", x"92119311", x"94119511", x"96119711",
		x"98119911", x"9A119B11", x"9C119D11", x"9E119F11", x"A011A111", x"A211A311", x"A411A511", x"A611A711",
		x"A811A911", x"AA11AB11", x"AC11AD11", x"AE11AF11", x"B011B111", x"B211B311", x"B411B511", x"B611B711",
		x"B811B911", x"BA11BB11", x"BC11BD11", x"BE11BF11", x"FFFFFFFF", x"FFFFFFFF", x"C011C111", x"C211C311",
		x"C411C511", x"C611C711", x"C811C911", x"CA11CB11", x"CC11CD11", x"CE11CF11", x"D011D111", x"D211D311",
		x"D411D511", x"D611D711", x"D811D911", x"DA11DB11", x"DC11DD11", x"DE11DF11", x"E011E111", x"E211E311",
		x"E411E511", x"E611E711", x"E811E911", x"EA11EB11", x"EC11ED11", x"EE11EF11", x"F011F111", x"F211F311",
		x"F411F511", x"F611F711", x"F811F911", x"FA11FB11", x"FC11FD11", x"FE11FF11", x"FFFFFFFF", x"FFFFFFFF",
		x"00120112", x"02120312", x"04120512", x"06120712", x"08120912", x"0A120B12", x"0C120D12", x"0E120F12",
		x"10121112", x"12121312", x"14121512", x"16121712", x"18121912", x"1A121B12", x"1C121D12", x"1E121F12",
		x"20122112", x"22122312", x"24122512", x"26122712", x"28122912", x"2A122B12", x"2C122D12", x"2E122F12",
		x"30123112", x"32123312", x"34123512", x"36123712", x"38123912", x"3A123B12", x"3C123D12", x"3E123F12",
		x"FFFFFFFF", x"FFFFFFFF", x"40124112", x"42124312", x"44124512", x"46124712", x"48124912", x"4A124B12",
		x"4C124D12", x"4E124F12", x"50125112", x"52125312", x"54125512", x"56125712", x"58125912", x"5A125B12",
		x"5C125D12", x"5E125F12", x"60126112", x"62126312", x"64126512", x"66126712", x"68126912", x"6A126B12",
		x"6C126D12", x"6E126F12", x"70127112", x"72127312", x"74127512", x"76127712", x"78127912", x"7A127B12",
		x"7C127D12", x"7E127F12", x"FFFFFFFF", x"FFFFFFFF", x"80128112", x"82128312", x"84128512", x"86128712",
		x"88128912", x"8A128B12", x"8C128D12", x"8E128F12", x"90129112", x"92129312", x"94129512", x"96129712",
		x"98129912", x"9A129B12", x"9C129D12", x"9E129F12", x"A012A112", x"A212A312", x"A412A512", x"A612A712",
		x"A812A912", x"AA12AB12", x"AC12AD12", x"AE12AF12", x"B012B112", x"B212B312", x"B412B512", x"B612B712",
		x"B812B912", x"BA12BB12", x"BC12BD12", x"BE12BF12", x"FFFFFFFF", x"FFFFFFFF", x"C012C112", x"C212C312",
		x"C412C512", x"C612C712", x"C812C912", x"CA12CB12", x"CC12CD12", x"CE12CF12", x"D012D112", x"D212D312",
		x"D412D512", x"D612D712", x"D812D912", x"DA12DB12", x"DC12DD12", x"DE12DF12", x"E012E112", x"E212E312",
		x"E412E512", x"E612E712", x"E812E912", x"EA12EB12", x"EC12ED12", x"EE12EF12", x"F012F112", x"F212F312",
		x"F412F512", x"F612F712", x"F812F912", x"FA12FB12", x"FC12FD12", x"FE12FF12", x"FFFFFFFF", x"FFFFFFFF",
		x"00130113", x"02130313", x"04130513", x"06130713", x"08130913", x"0A130B13", x"0C130D13", x"0E130F13",
		x"10131113", x"12131313", x"14131513", x"16131713", x"18131913", x"1A131B13", x"1C131D13", x"1E131F13",
		x"20132113", x"22132313", x"24132513", x"26132713", x"28132913", x"2A132B13", x"2C132D13", x"2E132F13",
		x"30133113", x"32133313", x"34133513", x"36133713", x"38133913", x"3A133B13", x"3C133D13", x"3E133F13",
		x"FFFFFFFF", x"FFFFFFFF", x"40134113", x"42134313", x"44134513", x"46134713", x"48134913", x"4A134B13",
		x"4C134D13", x"4E134F13", x"50135113", x"52135313", x"54135513", x"56135713", x"58135913", x"5A135B13",
		x"5C135D13", x"5E135F13", x"60136113", x"62136313", x"64136513", x"66136713", x"68136913", x"6A136B13",
		x"6C136D13", x"6E136F13", x"70137113", x"72137313", x"74137513", x"76137713", x"78137913", x"7A137B13",
		x"7C137D13", x"7E137F13", x"FFFFFFFF", x"FFFFFFFF", x"80138113", x"82138313", x"84138513", x"86138713",
		x"88138913", x"8A138B13", x"8C138D13", x"8E138F13", x"90139113", x"92139313", x"94139513", x"96139713",
		x"98139913", x"9A139B13", x"9C139D13", x"9E139F13", x"A013A113", x"A213A313", x"A413A513", x"A613A713",
		x"A813A913", x"AA13AB13", x"AC13AD13", x"AE13AF13", x"B013B113", x"B213B313", x"B413B513", x"B613B713",
		x"B813B913", x"BA13BB13", x"BC13BD13", x"BE13BF13", x"FFFFFFFF", x"FFFFFFFF", x"C013C113", x"C213C313",
		x"C413C513", x"C613C713", x"C813C913", x"CA13CB13", x"CC13CD13", x"CE13CF13", x"D013D113", x"D213D313",
		x"D413D513", x"D613D713", x"D813D913", x"DA13DB13", x"DC13DD13", x"DE13DF13", x"E013E113", x"E213E313",
		x"E413E513", x"E613E713", x"E813E913", x"EA13EB13", x"EC13ED13", x"EE13EF13", x"F013F113", x"F213F313",
		x"F413F513", x"F613F713", x"F813F913", x"FA13FB13", x"FC13FD13", x"FE13FF13", x"FFFFFFFF", x"FFFFFFFF",
		x"00140114", x"02140314", x"04140514", x"06140714", x"08140914", x"0A140B14", x"0C140D14", x"0E140F14",
		x"10141114", x"12141314", x"14141514", x"16141714", x"18141914", x"1A141B14", x"1C141D14", x"1E141F14",
		x"20142114", x"22142314", x"24142514", x"26142714", x"28142914", x"2A142B14", x"2C142D14", x"2E142F14",
		x"30143114", x"32143314", x"34143514", x"36143714", x"38143914", x"3A143B14", x"3C143D14", x"3E143F14",
		x"FFFFFFFF", x"FFFFFFFF", x"40144114", x"42144314", x"44144514", x"46144714", x"48144914", x"4A144B14",
		x"4C144D14", x"4E144F14", x"50145114", x"52145314", x"54145514", x"56145714", x"58145914", x"5A145B14",
		x"5C145D14", x"5E145F14", x"60146114", x"62146314", x"64146514", x"66146714", x"68146914", x"6A146B14",
		x"6C146D14", x"6E146F14", x"70147114", x"72147314", x"74147514", x"76147714", x"78147914", x"7A147B14",
		x"7C147D14", x"7E147F14", x"FFFFFFFF", x"FFFFFFFF", x"80148114", x"82148314", x"84148514", x"86148714",
		x"88148914", x"8A148B14", x"8C148D14", x"8E148F14", x"90149114", x"92149314", x"94149514", x"96149714",
		x"98149914", x"9A149B14", x"9C149D14", x"9E149F14", x"A014A114", x"A214A314", x"A414A514", x"A614A714",
		x"A814A914", x"AA14AB14", x"AC14AD14", x"AE14AF14", x"B014B114", x"B214B314", x"B414B514", x"B614B714",
		x"B814B914", x"BA14BB14", x"BC14BD14", x"BE14BF14", x"FFFFFFFF", x"FFFFFFFF", x"C014C114", x"C214C314",
		x"C414C514", x"C614C714", x"C814C914", x"CA14CB14", x"CC14CD14", x"CE14CF14", x"D014D114", x"D214D314",
		x"D414D514", x"D614D714", x"D814D914", x"DA14DB14", x"DC14DD14", x"DE14DF14", x"E014E114", x"E214E314",
		x"E414E514", x"E614E714", x"E814E914", x"EA14EB14", x"EC14ED14", x"EE14EF14", x"F014F114", x"F214F314",
		x"F414F514", x"F614F714", x"F814F914", x"FA14FB14", x"FC14FD14", x"FE14FF14", x"FFFFFFFF", x"FFFFFFFF",
		x"00150115", x"02150315", x"04150515", x"06150715", x"08150915", x"0A150B15", x"0C150D15", x"0E150F15",
		x"10151115", x"12151315", x"14151515", x"16151715", x"18151915", x"1A151B15", x"1C151D15", x"1E151F15",
		x"20152115", x"22152315", x"24152515", x"26152715", x"28152915", x"2A152B15", x"2C152D15", x"2E152F15",
		x"30153115", x"32153315", x"34153515", x"36153715", x"38153915", x"3A153B15", x"3C153D15", x"3E153F15",
		x"FFFFFFFF", x"FFFFFFFF", x"40154115", x"42154315", x"44154515", x"46154715", x"48154915", x"4A154B15",
		x"4C154D15", x"4E154F15", x"50155115", x"52155315", x"54155515", x"56155715", x"58155915", x"5A155B15",
		x"5C155D15", x"5E155F15", x"60156115", x"62156315", x"64156515", x"66156715", x"68156915", x"6A156B15",
		x"6C156D15", x"6E156F15", x"70157115", x"72157315", x"74157515", x"76157715", x"78157915", x"7A157B15",
		x"7C157D15", x"7E157F15", x"FFFFFFFF", x"FFFFFFFF", x"80158115", x"82158315", x"84158515", x"86158715",
		x"88158915", x"8A158B15", x"8C158D15", x"8E158F15", x"90159115", x"92159315", x"94159515", x"96159715",
		x"98159915", x"9A159B15", x"9C159D15", x"9E159F15", x"A015A115", x"A215A315", x"A415A515", x"A615A715",
		x"A815A915", x"AA15AB15", x"AC15AD15", x"AE15AF15", x"B015B115", x"B215B315", x"B415B515", x"B615B715",
		x"B815B915", x"BA15BB15", x"BC15BD15", x"BE15BF15", x"FFFFFFFF", x"FFFFFFFF", x"C015C115", x"C215C315",
		x"C415C515", x"C615C715", x"C815C915", x"CA15CB15", x"CC15CD15", x"CE15CF15", x"D015D115", x"D215D315",
		x"D415D515", x"D615D715", x"D815D915", x"DA15DB15", x"DC15DD15", x"DE15DF15", x"E015E115", x"E215E315",
		x"E415E515", x"E615E715", x"E815E915", x"EA15EB15", x"EC15ED15", x"EE15EF15", x"F015F115", x"F215F315",
		x"F415F515", x"F615F715", x"F815F915", x"FA15FB15", x"FC15FD15", x"FE15FF15", x"FFFFFFFF", x"FFFFFFFF",
		x"00160116", x"02160316", x"04160516", x"06160716", x"08160916", x"0A160B16", x"0C160D16", x"0E160F16",
		x"10161116", x"12161316", x"14161516", x"16161716", x"18161916", x"1A161B16", x"1C161D16", x"1E161F16",
		x"20162116", x"22162316", x"24162516", x"26162716", x"28162916", x"2A162B16", x"2C162D16", x"2E162F16",
		x"30163116", x"32163316", x"34163516", x"36163716", x"38163916", x"3A163B16", x"3C163D16", x"3E163F16",
		x"FFFFFFFF", x"FFFFFFFF", x"40164116", x"42164316", x"44164516", x"46164716", x"48164916", x"4A164B16",
		x"4C164D16", x"4E164F16", x"50165116", x"52165316", x"54165516", x"56165716", x"58165916", x"5A165B16",
		x"5C165D16", x"5E165F16", x"60166116", x"62166316", x"64166516", x"66166716", x"68166916", x"6A166B16",
		x"6C166D16", x"6E166F16", x"70167116", x"72167316", x"74167516", x"76167716", x"78167916", x"7A167B16",
		x"7C167D16", x"7E167F16", x"FFFFFFFF", x"FFFFFFFF", x"80168116", x"82168316", x"84168516", x"86168716",
		x"88168916", x"8A168B16", x"8C168D16", x"8E168F16", x"90169116", x"92169316", x"94169516", x"96169716",
		x"98169916", x"9A169B16", x"9C169D16", x"9E169F16", x"A016A116", x"A216A316", x"A416A516", x"A616A716",
		x"A816A916", x"AA16AB16", x"AC16AD16", x"AE16AF16", x"B016B116", x"B216B316", x"B416B516", x"B616B716",
		x"B816B916", x"BA16BB16", x"BC16BD16", x"BE16BF16", x"FFFFFFFF", x"FFFFFFFF", x"C016C116", x"C216C316",
		x"C416C516", x"C616C716", x"C816C916", x"CA16CB16", x"CC16CD16", x"CE16CF16", x"D016D116", x"D216D316",
		x"D416D516", x"D616D716", x"D816D916", x"DA16DB16", x"DC16DD16", x"DE16DF16", x"E016E116", x"E216E316",
		x"E416E516", x"E616E716", x"E816E916", x"EA16EB16", x"EC16ED16", x"EE16EF16", x"F016F116", x"F216F316",
		x"F416F516", x"F616F716", x"F816F916", x"FA16FB16", x"FC16FD16", x"FE16FF16", x"FFFFFFFF", x"FFFFFFFF",
		x"00170117", x"02170317", x"04170517", x"06170717", x"08170917", x"0A170B17", x"0C170D17", x"0E170F17",
		x"10171117", x"12171317", x"14171517", x"16171717", x"18171917", x"1A171B17", x"1C171D17", x"1E171F17",
		x"20172117", x"22172317", x"24172517", x"26172717", x"28172917", x"2A172B17", x"2C172D17", x"2E172F17",
		x"30173117", x"32173317", x"34173517", x"36173717", x"38173917", x"3A173B17", x"3C173D17", x"3E173F17",
		x"FFFFFFFF", x"FFFFFFFF", x"40174117", x"42174317", x"44174517", x"46174717", x"48174917", x"4A174B17",
		x"4C174D17", x"4E174F17", x"50175117", x"52175317", x"54175517", x"56175717", x"58175917", x"5A175B17",
		x"5C175D17", x"5E175F17", x"60176117", x"62176317", x"64176517", x"66176717", x"68176917", x"6A176B17",
		x"6C176D17", x"6E176F17", x"70177117", x"72177317", x"74177517", x"76177717", x"78177917", x"7A177B17",
		x"7C177D17", x"7E177F17", x"FFFFFFFF", x"FFFFFFFF", x"80178117", x"82178317", x"84178517", x"86178717",
		x"88178917", x"8A178B17", x"8C178D17", x"8E178F17", x"90179117", x"92179317", x"94179517", x"96179717",
		x"98179917", x"9A179B17", x"9C179D17", x"9E179F17", x"A017A117", x"A217A317", x"A417A517", x"A617A717",
		x"A817A917", x"AA17AB17", x"AC17AD17", x"AE17AF17", x"B017B117", x"B217B317", x"B417B517", x"B617B717",
		x"B817B917", x"BA17BB17", x"BC17BD17", x"BE17BF17", x"FFFFFFFF", x"FFFFFFFF", x"C017C117", x"C217C317",
		x"C417C517", x"C617C717", x"C817C917", x"CA17CB17", x"CC17CD17", x"CE17CF17", x"D017D117", x"D217D317",
		x"D417D517", x"D617D717", x"D817D917", x"DA17DB17", x"DC17DD17", x"DE17DF17", x"E017E117", x"E217E317",
		x"E417E517", x"E617E717", x"E817E917", x"EA17EB17", x"EC17ED17", x"EE17EF17", x"F017F117", x"F217F317",
		x"F417F517", x"F617F717", x"F817F917", x"FA17FB17", x"FC17FD17", x"FE17FF17", x"FFFFFFFF", x"FFFFFFFF",
		x"00180118", x"02180318", x"04180518", x"06180718", x"08180918", x"0A180B18", x"0C180D18", x"0E180F18",
		x"10181118", x"12181318", x"14181518", x"16181718", x"18181918", x"1A181B18", x"1C181D18", x"1E181F18",
		x"20182118", x"22182318", x"24182518", x"26182718", x"28182918", x"2A182B18", x"2C182D18", x"2E182F18",
		x"30183118", x"32183318", x"34183518", x"36183718", x"38183918", x"3A183B18", x"3C183D18", x"3E183F18",
		x"FFFFFFFF", x"FFFFFFFF", x"40184118", x"42184318", x"44184518", x"46184718", x"48184918", x"4A184B18",
		x"4C184D18", x"4E184F18", x"50185118", x"52185318", x"54185518", x"56185718", x"58185918", x"5A185B18",
		x"5C185D18", x"5E185F18", x"60186118", x"62186318", x"64186518", x"66186718", x"68186918", x"6A186B18",
		x"6C186D18", x"6E186F18", x"70187118", x"72187318", x"74187518", x"76187718", x"78187918", x"7A187B18",
		x"7C187D18", x"7E187F18", x"FFFFFFFF", x"FFFFFFFF", x"80188118", x"82188318", x"84188518", x"86188718",
		x"88188918", x"8A188B18", x"8C188D18", x"8E188F18", x"90189118", x"92189318", x"94189518", x"96189718",
		x"98189918", x"9A189B18", x"9C189D18", x"9E189F18", x"A018A118", x"A218A318", x"A418A518", x"A618A718",
		x"A818A918", x"AA18AB18", x"AC18AD18", x"AE18AF18", x"B018B118", x"B218B318", x"B418B518", x"B618B718",
		x"B818B918", x"BA18BB18", x"BC18BD18", x"BE18BF18", x"FFFFFFFF", x"FFFFFFFF", x"C018C118", x"C218C318",
		x"C418C518", x"C618C718", x"C818C918", x"CA18CB18", x"CC18CD18", x"CE18CF18", x"D018D118", x"D218D318",
		x"D418D518", x"D618D718", x"D818D918", x"DA18DB18", x"DC18DD18", x"DE18DF18", x"E018E118", x"E218E318",
		x"E418E518", x"E618E718", x"E818E918", x"EA18EB18", x"EC18ED18", x"EE18EF18", x"F018F118", x"F218F318",
		x"F418F518", x"F618F718", x"F818F918", x"FA18FB18", x"FC18FD18", x"FE18FF18", x"FFFFFFFF", x"FFFFFFFF",
		x"00190119", x"02190319", x"04190519", x"06190719", x"08190919", x"0A190B19", x"0C190D19", x"0E190F19",
		x"10191119", x"12191319", x"14191519", x"16191719", x"18191919", x"1A191B19", x"1C191D19", x"1E191F19",
		x"20192119", x"22192319", x"24192519", x"26192719", x"28192919", x"2A192B19", x"2C192D19", x"2E192F19",
		x"30193119", x"32193319", x"34193519", x"36193719", x"38193919", x"3A193B19", x"3C193D19", x"3E193F19",
		x"FFFFFFFF", x"FFFFFFFF", x"40194119", x"42194319", x"44194519", x"46194719", x"48194919", x"4A194B19",
		x"4C194D19", x"4E194F19", x"50195119", x"52195319", x"54195519", x"56195719", x"58195919", x"5A195B19",
		x"5C195D19", x"5E195F19", x"60196119", x"62196319", x"64196519", x"66196719", x"68196919", x"6A196B19",
		x"6C196D19", x"6E196F19", x"70197119", x"72197319", x"74197519", x"76197719", x"78197919", x"7A197B19",
		x"7C197D19", x"7E197F19", x"FFFFFFFF", x"FFFFFFFF", x"80198119", x"82198319", x"84198519", x"86198719",
		x"88198919", x"8A198B19", x"8C198D19", x"8E198F19", x"90199119", x"92199319", x"94199519", x"96199719",
		x"98199919", x"9A199B19", x"9C199D19", x"9E199F19", x"A019A119", x"A219A319", x"A419A519", x"A619A719",
		x"A819A919", x"AA19AB19", x"AC19AD19", x"AE19AF19", x"B019B119", x"B219B319", x"B419B519", x"B619B719",
		x"B819B919", x"BA19BB19", x"BC19BD19", x"BE19BF19", x"FFFFFFFF", x"FFFFFFFF", x"C019C119", x"C219C319",
		x"C419C519", x"C619C719", x"C819C919", x"CA19CB19", x"CC19CD19", x"CE19CF19", x"D019D119", x"D219D319",
		x"D419D519", x"D619D719", x"D819D919", x"DA19DB19", x"DC19DD19", x"DE19DF19", x"E019E119", x"E219E319",
		x"E419E519", x"E619E719", x"E819E919", x"EA19EB19", x"EC19ED19", x"EE19EF19", x"F019F119", x"F219F319",
		x"F419F519", x"F619F719", x"F819F919", x"FA19FB19", x"FC19FD19", x"FE19FF19", x"FFFFFFFF", x"FFFFFFFF",
		x"001A011A", x"021A031A", x"041A051A", x"061A071A", x"081A091A", x"0A1A0B1A", x"0C1A0D1A", x"0E1A0F1A",
		x"101A111A", x"121A131A", x"141A151A", x"161A171A", x"181A191A", x"1A1A1B1A", x"1C1A1D1A", x"1E1A1F1A",
		x"201A211A", x"221A231A", x"241A251A", x"261A271A", x"281A291A", x"2A1A2B1A", x"2C1A2D1A", x"2E1A2F1A",
		x"301A311A", x"321A331A", x"341A351A", x"361A371A", x"381A391A", x"3A1A3B1A", x"3C1A3D1A", x"3E1A3F1A",
		x"FFFFFFFF", x"FFFFFFFF", x"401A411A", x"421A431A", x"441A451A", x"461A471A", x"481A491A", x"4A1A4B1A",
		x"4C1A4D1A", x"4E1A4F1A", x"501A511A", x"521A531A", x"541A551A", x"561A571A", x"581A591A", x"5A1A5B1A",
		x"5C1A5D1A", x"5E1A5F1A", x"601A611A", x"621A631A", x"641A651A", x"661A671A", x"681A691A", x"6A1A6B1A",
		x"6C1A6D1A", x"6E1A6F1A", x"701A711A", x"721A731A", x"741A751A", x"761A771A", x"781A791A", x"7A1A7B1A",
		x"7C1A7D1A", x"7E1A7F1A", x"FFFFFFFF", x"FFFFFFFF", x"801A811A", x"821A831A", x"841A851A", x"861A871A",
		x"881A891A", x"8A1A8B1A", x"8C1A8D1A", x"8E1A8F1A", x"901A911A", x"921A931A", x"941A951A", x"961A971A",
		x"981A991A", x"9A1A9B1A", x"9C1A9D1A", x"9E1A9F1A", x"A01AA11A", x"A21AA31A", x"A41AA51A", x"A61AA71A",
		x"A81AA91A", x"AA1AAB1A", x"AC1AAD1A", x"AE1AAF1A", x"B01AB11A", x"B21AB31A", x"B41AB51A", x"B61AB71A",
		x"B81AB91A", x"BA1ABB1A", x"BC1ABD1A", x"BE1ABF1A", x"FFFFFFFF", x"FFFFFFFF", x"C01AC11A", x"C21AC31A",
		x"C41AC51A", x"C61AC71A", x"C81AC91A", x"CA1ACB1A", x"CC1ACD1A", x"CE1ACF1A", x"D01AD11A", x"D21AD31A",
		x"D41AD51A", x"D61AD71A", x"D81AD91A", x"DA1ADB1A", x"DC1ADD1A", x"DE1ADF1A", x"E01AE11A", x"E21AE31A",
		x"E41AE51A", x"E61AE71A", x"E81AE91A", x"EA1AEB1A", x"EC1AED1A", x"EE1AEF1A", x"F01AF11A", x"F21AF31A",
		x"F41AF51A", x"F61AF71A", x"F81AF91A", x"FA1AFB1A", x"FC1AFD1A", x"FE1AFF1A", x"FFFFFFFF", x"FFFFFFFF",
		x"001B011B", x"021B031B", x"041B051B", x"061B071B", x"081B091B", x"0A1B0B1B", x"0C1B0D1B", x"0E1B0F1B",
		x"101B111B", x"121B131B", x"141B151B", x"161B171B", x"181B191B", x"1A1B1B1B", x"1C1B1D1B", x"1E1B1F1B",
		x"201B211B", x"221B231B", x"241B251B", x"261B271B", x"281B291B", x"2A1B2B1B", x"2C1B2D1B", x"2E1B2F1B",
		x"301B311B", x"321B331B", x"341B351B", x"361B371B", x"381B391B", x"3A1B3B1B", x"3C1B3D1B", x"3E1B3F1B",
		x"FFFFFFFF", x"FFFFFFFF", x"401B411B", x"421B431B", x"441B451B", x"461B471B", x"481B491B", x"4A1B4B1B",
		x"4C1B4D1B", x"4E1B4F1B", x"501B511B", x"521B531B", x"541B551B", x"561B571B", x"581B591B", x"5A1B5B1B",
		x"5C1B5D1B", x"5E1B5F1B", x"601B611B", x"621B631B", x"641B651B", x"661B671B", x"681B691B", x"6A1B6B1B",
		x"6C1B6D1B", x"6E1B6F1B", x"701B711B", x"721B731B", x"741B751B", x"761B771B", x"781B791B", x"7A1B7B1B",
		x"7C1B7D1B", x"7E1B7F1B", x"FFFFFFFF", x"FFFFFFFF", x"801B811B", x"821B831B", x"841B851B", x"861B871B",
		x"881B891B", x"8A1B8B1B", x"8C1B8D1B", x"8E1B8F1B", x"901B911B", x"921B931B", x"941B951B", x"961B971B",
		x"981B991B", x"9A1B9B1B", x"9C1B9D1B", x"9E1B9F1B", x"A01BA11B", x"A21BA31B", x"A41BA51B", x"A61BA71B",
		x"A81BA91B", x"AA1BAB1B", x"AC1BAD1B", x"AE1BAF1B", x"B01BB11B", x"B21BB31B", x"B41BB51B", x"B61BB71B",
		x"B81BB91B", x"BA1BBB1B", x"BC1BBD1B", x"BE1BBF1B", x"FFFFFFFF", x"FFFFFFFF", x"C01BC11B", x"C21BC31B",
		x"C41BC51B", x"C61BC71B", x"C81BC91B", x"CA1BCB1B", x"CC1BCD1B", x"CE1BCF1B", x"D01BD11B", x"D21BD31B",
		x"D41BD51B", x"D61BD71B", x"D81BD91B", x"DA1BDB1B", x"DC1BDD1B", x"DE1BDF1B", x"E01BE11B", x"E21BE31B",
		x"E41BE51B", x"E61BE71B", x"E81BE91B", x"EA1BEB1B", x"EC1BED1B", x"EE1BEF1B", x"F01BF11B", x"F21BF31B",
		x"F41BF51B", x"F61BF71B", x"F81BF91B", x"FA1BFB1B", x"FC1BFD1B", x"FE1BFF1B", x"FFFFFFFF", x"FFFFFFFF",
		x"001C011C", x"021C031C", x"041C051C", x"061C071C", x"081C091C", x"0A1C0B1C", x"0C1C0D1C", x"0E1C0F1C",
		x"101C111C", x"121C131C", x"141C151C", x"161C171C", x"181C191C", x"1A1C1B1C", x"1C1C1D1C", x"1E1C1F1C",
		x"201C211C", x"221C231C", x"241C251C", x"261C271C", x"281C291C", x"2A1C2B1C", x"2C1C2D1C", x"2E1C2F1C",
		x"301C311C", x"321C331C", x"341C351C", x"361C371C", x"381C391C", x"3A1C3B1C", x"3C1C3D1C", x"3E1C3F1C",
		x"FFFFFFFF", x"FFFFFFFF", x"401C411C", x"421C431C", x"441C451C", x"461C471C", x"481C491C", x"4A1C4B1C",
		x"4C1C4D1C", x"4E1C4F1C", x"501C511C", x"521C531C", x"541C551C", x"561C571C", x"581C591C", x"5A1C5B1C",
		x"5C1C5D1C", x"5E1C5F1C", x"601C611C", x"621C631C", x"641C651C", x"661C671C", x"681C691C", x"6A1C6B1C",
		x"6C1C6D1C", x"6E1C6F1C", x"701C711C", x"721C731C", x"741C751C", x"761C771C", x"781C791C", x"7A1C7B1C",
		x"7C1C7D1C", x"7E1C7F1C", x"FFFFFFFF", x"FFFFFFFF", x"801C811C", x"821C831C", x"841C851C", x"861C871C",
		x"881C891C", x"8A1C8B1C", x"8C1C8D1C", x"8E1C8F1C", x"901C911C", x"921C931C", x"941C951C", x"961C971C",
		x"981C991C", x"9A1C9B1C", x"9C1C9D1C", x"9E1C9F1C", x"A01CA11C", x"A21CA31C", x"A41CA51C", x"A61CA71C",
		x"A81CA91C", x"AA1CAB1C", x"AC1CAD1C", x"AE1CAF1C", x"B01CB11C", x"B21CB31C", x"B41CB51C", x"B61CB71C",
		x"B81CB91C", x"BA1CBB1C", x"BC1CBD1C", x"BE1CBF1C", x"FFFFFFFF", x"FFFFFFFF", x"C01CC11C", x"C21CC31C",
		x"C41CC51C", x"C61CC71C", x"C81CC91C", x"CA1CCB1C", x"CC1CCD1C", x"CE1CCF1C", x"D01CD11C", x"D21CD31C",
		x"D41CD51C", x"D61CD71C", x"D81CD91C", x"DA1CDB1C", x"DC1CDD1C", x"DE1CDF1C", x"E01CE11C", x"E21CE31C",
		x"E41CE51C", x"E61CE71C", x"E81CE91C", x"EA1CEB1C", x"EC1CED1C", x"EE1CEF1C", x"F01CF11C", x"F21CF31C",
		x"F41CF51C", x"F61CF71C", x"F81CF91C", x"FA1CFB1C", x"FC1CFD1C", x"FE1CFF1C", x"FFFFFFFF", x"FFFFFFFF",
		x"001D011D", x"021D031D", x"041D051D", x"061D071D", x"081D091D", x"0A1D0B1D", x"0C1D0D1D", x"0E1D0F1D",
		x"101D111D", x"121D131D", x"141D151D", x"161D171D", x"181D191D", x"1A1D1B1D", x"1C1D1D1D", x"1E1D1F1D",
		x"201D211D", x"221D231D", x"241D251D", x"261D271D", x"281D291D", x"2A1D2B1D", x"2C1D2D1D", x"2E1D2F1D",
		x"301D311D", x"321D331D", x"341D351D", x"361D371D", x"381D391D", x"3A1D3B1D", x"3C1D3D1D", x"3E1D3F1D",
		x"FFFFFFFF", x"FFFFFFFF", x"401D411D", x"421D431D", x"441D451D", x"461D471D", x"481D491D", x"4A1D4B1D",
		x"4C1D4D1D", x"4E1D4F1D", x"501D511D", x"521D531D", x"541D551D", x"561D571D", x"581D591D", x"5A1D5B1D",
		x"5C1D5D1D", x"5E1D5F1D", x"601D611D", x"621D631D", x"641D651D", x"661D671D", x"681D691D", x"6A1D6B1D",
		x"6C1D6D1D", x"6E1D6F1D", x"701D711D", x"721D731D", x"741D751D", x"761D771D", x"781D791D", x"7A1D7B1D",
		x"7C1D7D1D", x"7E1D7F1D", x"FFFFFFFF", x"FFFFFFFF", x"801D811D", x"821D831D", x"841D851D", x"861D871D",
		x"881D891D", x"8A1D8B1D", x"8C1D8D1D", x"8E1D8F1D", x"901D911D", x"921D931D", x"941D951D", x"961D971D",
		x"981D991D", x"9A1D9B1D", x"9C1D9D1D", x"9E1D9F1D", x"A01DA11D", x"A21DA31D", x"A41DA51D", x"A61DA71D",
		x"A81DA91D", x"AA1DAB1D", x"AC1DAD1D", x"AE1DAF1D", x"B01DB11D", x"B21DB31D", x"B41DB51D", x"B61DB71D",
		x"B81DB91D", x"BA1DBB1D", x"BC1DBD1D", x"BE1DBF1D", x"FFFFFFFF", x"FFFFFFFF", x"C01DC11D", x"C21DC31D",
		x"C41DC51D", x"C61DC71D", x"C81DC91D", x"CA1DCB1D", x"CC1DCD1D", x"CE1DCF1D", x"D01DD11D", x"D21DD31D",
		x"D41DD51D", x"D61DD71D", x"D81DD91D", x"DA1DDB1D", x"DC1DDD1D", x"DE1DDF1D", x"E01DE11D", x"E21DE31D",
		x"E41DE51D", x"E61DE71D", x"E81DE91D", x"EA1DEB1D", x"EC1DED1D", x"EE1DEF1D", x"F01DF11D", x"F21DF31D",
		x"F41DF51D", x"F61DF71D", x"F81DF91D", x"FA1DFB1D", x"FC1DFD1D", x"FE1DFF1D", x"FFFFFFFF", x"FFFFFFFF",
		x"001E011E", x"021E031E", x"041E051E", x"061E071E", x"081E091E", x"0A1E0B1E", x"0C1E0D1E", x"0E1E0F1E",
		x"101E111E", x"121E131E", x"141E151E", x"161E171E", x"181E191E", x"1A1E1B1E", x"1C1E1D1E", x"1E1E1F1E",
		x"201E211E", x"221E231E", x"241E251E", x"261E271E", x"281E291E", x"2A1E2B1E", x"2C1E2D1E", x"2E1E2F1E",
		x"301E311E", x"321E331E", x"341E351E", x"361E371E", x"381E391E", x"3A1E3B1E", x"3C1E3D1E", x"3E1E3F1E",
		x"FFFFFFFF", x"FFFFFFFF", x"401E411E", x"421E431E", x"441E451E", x"461E471E", x"481E491E", x"4A1E4B1E",
		x"4C1E4D1E", x"4E1E4F1E", x"501E511E", x"521E531E", x"541E551E", x"561E571E", x"581E591E", x"5A1E5B1E",
		x"5C1E5D1E", x"5E1E5F1E", x"601E611E", x"621E631E", x"641E651E", x"661E671E", x"681E691E", x"6A1E6B1E",
		x"6C1E6D1E", x"6E1E6F1E", x"701E711E", x"721E731E", x"741E751E", x"761E771E", x"781E791E", x"7A1E7B1E",
		x"7C1E7D1E", x"7E1E7F1E", x"FFFFFFFF", x"FFFFFFFF", x"801E811E", x"821E831E", x"841E851E", x"861E871E",
		x"881E891E", x"8A1E8B1E", x"8C1E8D1E", x"8E1E8F1E", x"901E911E", x"921E931E", x"941E951E", x"961E971E",
		x"981E991E", x"9A1E9B1E", x"9C1E9D1E", x"9E1E9F1E", x"A01EA11E", x"A21EA31E", x"A41EA51E", x"A61EA71E",
		x"A81EA91E", x"AA1EAB1E", x"AC1EAD1E", x"AE1EAF1E", x"B01EB11E", x"B21EB31E", x"B41EB51E", x"B61EB71E",
		x"B81EB91E", x"BA1EBB1E", x"BC1EBD1E", x"BE1EBF1E", x"FFFFFFFF", x"FFFFFFFF", x"C01EC11E", x"C21EC31E",
		x"C41EC51E", x"C61EC71E", x"C81EC91E", x"CA1ECB1E", x"CC1ECD1E", x"CE1ECF1E", x"D01ED11E", x"D21ED31E",
		x"D41ED51E", x"D61ED71E", x"D81ED91E", x"DA1EDB1E", x"DC1EDD1E", x"DE1EDF1E", x"E01EE11E", x"E21EE31E",
		x"E41EE51E", x"E61EE71E", x"E81EE91E", x"EA1EEB1E", x"EC1EED1E", x"EE1EEF1E", x"F01EF11E", x"F21EF31E",
		x"F41EF51E", x"F61EF71E", x"F81EF91E", x"FA1EFB1E", x"FC1EFD1E", x"FE1EFF1E", x"FFFFFFFF", x"FFFFFFFF",
		x"001F011F", x"021F031F", x"041F051F", x"061F071F", x"081F091F", x"0A1F0B1F", x"0C1F0D1F", x"0E1F0F1F",
		x"101F111F", x"121F131F", x"141F151F", x"161F171F", x"181F191F", x"1A1F1B1F", x"1C1F1D1F", x"1E1F1F1F",
		x"201F211F", x"221F231F", x"241F251F", x"261F271F", x"281F291F", x"2A1F2B1F", x"2C1F2D1F", x"2E1F2F1F",
		x"301F311F", x"321F331F", x"341F351F", x"361F371F", x"381F391F", x"3A1F3B1F", x"3C1F3D1F", x"3E1F3F1F",
		x"FFFFFFFF", x"FFFFFFFF", x"401F411F", x"421F431F", x"441F451F", x"461F471F", x"481F491F", x"4A1F4B1F",
		x"4C1F4D1F", x"4E1F4F1F", x"501F511F", x"521F531F", x"541F551F", x"561F571F", x"581F591F", x"5A1F5B1F",
		x"5C1F5D1F", x"5E1F5F1F", x"601F611F", x"621F631F", x"641F651F", x"661F671F", x"681F691F", x"6A1F6B1F",
		x"6C1F6D1F", x"6E1F6F1F", x"701F711F", x"721F731F", x"741F751F", x"761F771F", x"781F791F", x"7A1F7B1F",
		x"7C1F7D1F", x"7E1F7F1F", x"FFFFFFFF", x"FFFFFFFF", x"801F811F", x"821F831F", x"841F851F", x"861F871F",
		x"881F891F", x"8A1F8B1F", x"8C1F8D1F", x"8E1F8F1F", x"901F911F", x"921F931F", x"941F951F", x"961F971F",
		x"981F991F", x"9A1F9B1F", x"9C1F9D1F", x"9E1F9F1F", x"A01FA11F", x"A21FA31F", x"A41FA51F", x"A61FA71F",
		x"A81FA91F", x"AA1FAB1F", x"AC1FAD1F", x"AE1FAF1F", x"B01FB11F", x"B21FB31F", x"B41FB51F", x"B61FB71F",
		x"B81FB91F", x"BA1FBB1F", x"BC1FBD1F", x"BE1FBF1F", x"FFFFFFFF", x"FFFFFFFF", x"C01FC11F", x"C21FC31F",
		x"C41FC51F", x"C61FC71F", x"C81FC91F", x"CA1FCB1F", x"CC1FCD1F", x"CE1FCF1F", x"D01FD11F", x"D21FD31F",
		x"D41FD51F", x"D61FD71F", x"D81FD91F", x"DA1FDB1F", x"DC1FDD1F", x"DE1FDF1F", x"E01FE11F", x"E21FE31F",
		x"E41FE51F", x"E61FE71F", x"E81FE91F", x"EA1FEB1F", x"EC1FED1F", x"EE1FEF1F", x"F01FF11F", x"F21FF31F",
		x"F41FF51F", x"F61FF71F", x"F81FF91F", x"FA1FFB1F", x"FC1FFD1F", x"FE1FFF1F", x"FFFFFFFF", x"FFFFFFFF",
		x"00200120", x"02200320", x"04200520", x"06200720", x"08200920", x"0A200B20", x"0C200D20", x"0E200F20",
		x"10201120", x"12201320", x"14201520", x"16201720", x"18201920", x"1A201B20", x"1C201D20", x"1E201F20",
		x"20202120", x"22202320", x"24202520", x"26202720", x"28202920", x"2A202B20", x"2C202D20", x"2E202F20",
		x"30203120", x"32203320", x"34203520", x"36203720", x"38203920", x"3A203B20", x"3C203D20", x"3E203F20",
		x"FFFFFFFF", x"FFFFFFFF", x"40204120", x"42204320", x"44204520", x"46204720", x"48204920", x"4A204B20",
		x"4C204D20", x"4E204F20", x"50205120", x"52205320", x"54205520", x"56205720", x"58205920", x"5A205B20",
		x"5C205D20", x"5E205F20", x"60206120", x"62206320", x"64206520", x"66206720", x"68206920", x"6A206B20",
		x"6C206D20", x"6E206F20", x"70207120", x"72207320", x"74207520", x"76207720", x"78207920", x"7A207B20",
		x"7C207D20", x"7E207F20", x"FFFFFFFF", x"FFFFFFFF", x"80208120", x"82208320", x"84208520", x"86208720",
		x"88208920", x"8A208B20", x"8C208D20", x"8E208F20", x"90209120", x"92209320", x"94209520", x"96209720",
		x"98209920", x"9A209B20", x"9C209D20", x"9E209F20", x"A020A120", x"A220A320", x"A420A520", x"A620A720",
		x"A820A920", x"AA20AB20", x"AC20AD20", x"AE20AF20", x"B020B120", x"B220B320", x"B420B520", x"B620B720",
		x"B820B920", x"BA20BB20", x"BC20BD20", x"BE20BF20", x"FFFFFFFF", x"FFFFFFFF", x"C020C120", x"C220C320",
		x"C420C520", x"C620C720", x"C820C920", x"CA20CB20", x"CC20CD20", x"CE20CF20", x"D020D120", x"D220D320",
		x"D420D520", x"D620D720", x"D820D920", x"DA20DB20", x"DC20DD20", x"DE20DF20", x"E020E120", x"E220E320",
		x"E420E520", x"E620E720", x"E820E920", x"EA20EB20", x"EC20ED20", x"EE20EF20", x"F020F120", x"F220F320",
		x"F420F520", x"F620F720", x"F820F920", x"FA20FB20", x"FC20FD20", x"FE20FF20", x"FFFFFFFF", x"FFFFFFFF",
		x"00210121", x"02210321", x"04210521", x"06210721", x"08210921", x"0A210B21", x"0C210D21", x"0E210F21",
		x"10211121", x"12211321", x"14211521", x"16211721", x"18211921", x"1A211B21", x"1C211D21", x"1E211F21",
		x"20212121", x"22212321", x"24212521", x"26212721", x"28212921", x"2A212B21", x"2C212D21", x"2E212F21",
		x"30213121", x"32213321", x"34213521", x"36213721", x"38213921", x"3A213B21", x"3C213D21", x"3E213F21",
		x"FFFFFFFF", x"FFFFFFFF", x"40214121", x"42214321", x"44214521", x"46214721", x"48214921", x"4A214B21",
		x"4C214D21", x"4E214F21", x"50215121", x"52215321", x"54215521", x"56215721", x"58215921", x"5A215B21",
		x"5C215D21", x"5E215F21", x"60216121", x"62216321", x"64216521", x"66216721", x"68216921", x"6A216B21",
		x"6C216D21", x"6E216F21", x"70217121", x"72217321", x"74217521", x"76217721", x"78217921", x"7A217B21",
		x"7C217D21", x"7E217F21", x"FFFFFFFF", x"FFFFFFFF", x"80218121", x"82218321", x"84218521", x"86218721",
		x"88218921", x"8A218B21", x"8C218D21", x"8E218F21", x"90219121", x"92219321", x"94219521", x"96219721",
		x"98219921", x"9A219B21", x"9C219D21", x"9E219F21", x"A021A121", x"A221A321", x"A421A521", x"A621A721",
		x"A821A921", x"AA21AB21", x"AC21AD21", x"AE21AF21", x"B021B121", x"B221B321", x"B421B521", x"B621B721",
		x"B821B921", x"BA21BB21", x"BC21BD21", x"BE21BF21", x"FFFFFFFF", x"FFFFFFFF", x"C021C121", x"C221C321",
		x"C421C521", x"C621C721", x"C821C921", x"CA21CB21", x"CC21CD21", x"CE21CF21", x"D021D121", x"D221D321",
		x"D421D521", x"D621D721", x"D821D921", x"DA21DB21", x"DC21DD21", x"DE21DF21", x"E021E121", x"E221E321",
		x"E421E521", x"E621E721", x"E821E921", x"EA21EB21", x"EC21ED21", x"EE21EF21", x"F021F121", x"F221F321",
		x"F421F521", x"F621F721", x"F821F921", x"FA21FB21", x"FC21FD21", x"FE21FF21", x"FFFFFFFF", x"FFFFFFFF",
		x"00220122", x"02220322", x"04220522", x"06220722", x"08220922", x"0A220B22", x"0C220D22", x"0E220F22",
		x"10221122", x"12221322", x"14221522", x"16221722", x"18221922", x"1A221B22", x"1C221D22", x"1E221F22",
		x"20222122", x"22222322", x"24222522", x"26222722", x"28222922", x"2A222B22", x"2C222D22", x"2E222F22",
		x"30223122", x"32223322", x"34223522", x"36223722", x"38223922", x"3A223B22", x"3C223D22", x"3E223F22",
		x"FFFFFFFF", x"FFFFFFFF", x"40224122", x"42224322", x"44224522", x"46224722", x"48224922", x"4A224B22",
		x"4C224D22", x"4E224F22", x"50225122", x"52225322", x"54225522", x"56225722", x"58225922", x"5A225B22",
		x"5C225D22", x"5E225F22", x"60226122", x"62226322", x"64226522", x"66226722", x"68226922", x"6A226B22",
		x"6C226D22", x"6E226F22", x"70227122", x"72227322", x"74227522", x"76227722", x"78227922", x"7A227B22",
		x"7C227D22", x"7E227F22", x"FFFFFFFF", x"FFFFFFFF", x"80228122", x"82228322", x"84228522", x"86228722",
		x"88228922", x"8A228B22", x"8C228D22", x"8E228F22", x"90229122", x"92229322", x"94229522", x"96229722",
		x"98229922", x"9A229B22", x"9C229D22", x"9E229F22", x"A022A122", x"A222A322", x"A422A522", x"A622A722",
		x"A822A922", x"AA22AB22", x"AC22AD22", x"AE22AF22", x"B022B122", x"B222B322", x"B422B522", x"B622B722",
		x"B822B922", x"BA22BB22", x"BC22BD22", x"BE22BF22", x"FFFFFFFF", x"FFFFFFFF", x"C022C122", x"C222C322",
		x"C422C522", x"C622C722", x"C822C922", x"CA22CB22", x"CC22CD22", x"CE22CF22", x"D022D122", x"D222D322",
		x"D422D522", x"D622D722", x"D822D922", x"DA22DB22", x"DC22DD22", x"DE22DF22", x"E022E122", x"E222E322",
		x"E422E522", x"E622E722", x"E822E922", x"EA22EB22", x"EC22ED22", x"EE22EF22", x"F022F122", x"F222F322",
		x"F422F522", x"F622F722", x"F822F922", x"FA22FB22", x"FC22FD22", x"FE22FF22", x"FFFFFFFF", x"FFFFFFFF",
		x"00230123", x"02230323", x"04230523", x"06230723", x"08230923", x"0A230B23", x"0C230D23", x"0E230F23",
		x"10231123", x"12231323", x"14231523", x"16231723", x"18231923", x"1A231B23", x"1C231D23", x"1E231F23",
		x"20232123", x"22232323", x"24232523", x"26232723", x"28232923", x"2A232B23", x"2C232D23", x"2E232F23",
		x"30233123", x"32233323", x"34233523", x"36233723", x"38233923", x"3A233B23", x"3C233D23", x"3E233F23",
		x"FFFFFFFF", x"FFFFFFFF", x"40234123", x"42234323", x"44234523", x"46234723", x"48234923", x"4A234B23",
		x"4C234D23", x"4E234F23", x"50235123", x"52235323", x"54235523", x"56235723", x"58235923", x"5A235B23",
		x"5C235D23", x"5E235F23", x"60236123", x"62236323", x"64236523", x"66236723", x"68236923", x"6A236B23",
		x"6C236D23", x"6E236F23", x"70237123", x"72237323", x"74237523", x"76237723", x"78237923", x"7A237B23",
		x"7C237D23", x"7E237F23", x"FFFFFFFF", x"FFFFFFFF", x"80238123", x"82238323", x"84238523", x"86238723",
		x"88238923", x"8A238B23", x"8C238D23", x"8E238F23", x"90239123", x"92239323", x"94239523", x"96239723",
		x"98239923", x"9A239B23", x"9C239D23", x"9E239F23", x"A023A123", x"A223A323", x"A423A523", x"A623A723",
		x"A823A923", x"AA23AB23", x"AC23AD23", x"AE23AF23", x"B023B123", x"B223B323", x"B423B523", x"B623B723",
		x"B823B923", x"BA23BB23", x"BC23BD23", x"BE23BF23", x"FFFFFFFF", x"FFFFFFFF", x"C023C123", x"C223C323",
		x"C423C523", x"C623C723", x"C823C923", x"CA23CB23", x"CC23CD23", x"CE23CF23", x"D023D123", x"D223D323",
		x"D423D523", x"D623D723", x"D823D923", x"DA23DB23", x"DC23DD23", x"DE23DF23", x"E023E123", x"E223E323",
		x"E423E523", x"E623E723", x"E823E923", x"EA23EB23", x"EC23ED23", x"EE23EF23", x"F023F123", x"F223F323",
		x"F423F523", x"F623F723", x"F823F923", x"FA23FB23", x"FC23FD23", x"FE23FF23", x"FFFFFFFF", x"FFFFFFFF",
		x"00240124", x"02240324", x"04240524", x"06240724", x"08240924", x"0A240B24", x"0C240D24", x"0E240F24",
		x"10241124", x"12241324", x"14241524", x"16241724", x"18241924", x"1A241B24", x"1C241D24", x"1E241F24",
		x"20242124", x"22242324", x"24242524", x"26242724", x"28242924", x"2A242B24", x"2C242D24", x"2E242F24",
		x"30243124", x"32243324", x"34243524", x"36243724", x"38243924", x"3A243B24", x"3C243D24", x"3E243F24",
		x"FFFFFFFF", x"FFFFFFFF", x"40244124", x"42244324", x"44244524", x"46244724", x"48244924", x"4A244B24",
		x"4C244D24", x"4E244F24", x"50245124", x"52245324", x"54245524", x"56245724", x"58245924", x"5A245B24",
		x"5C245D24", x"5E245F24", x"60246124", x"62246324", x"64246524", x"66246724", x"68246924", x"6A246B24",
		x"6C246D24", x"6E246F24", x"70247124", x"72247324", x"74247524", x"76247724", x"78247924", x"7A247B24",
		x"7C247D24", x"7E247F24", x"FFFFFFFF", x"FFFFFFFF", x"80248124", x"82248324", x"84248524", x"86248724",
		x"88248924", x"8A248B24", x"8C248D24", x"8E248F24", x"90249124", x"92249324", x"94249524", x"96249724",
		x"98249924", x"9A249B24", x"9C249D24", x"9E249F24", x"A024A124", x"A224A324", x"A424A524", x"A624A724",
		x"A824A924", x"AA24AB24", x"AC24AD24", x"AE24AF24", x"B024B124", x"B224B324", x"B424B524", x"B624B724",
		x"B824B924", x"BA24BB24", x"BC24BD24", x"BE24BF24", x"FFFFFFFF", x"FFFFFFFF", x"C024C124", x"C224C324",
		x"C424C524", x"C624C724", x"C824C924", x"CA24CB24", x"CC24CD24", x"CE24CF24", x"D024D124", x"D224D324",
		x"D424D524", x"D624D724", x"D824D924", x"DA24DB24", x"DC24DD24", x"DE24DF24", x"E024E124", x"E224E324",
		x"E424E524", x"E624E724", x"E824E924", x"EA24EB24", x"EC24ED24", x"EE24EF24", x"F024F124", x"F224F324",
		x"F424F524", x"F624F724", x"F824F924", x"FA24FB24", x"FC24FD24", x"FE24FF24", x"FFFFFFFF", x"FFFFFFFF",
		x"00250125", x"02250325", x"04250525", x"06250725", x"08250925", x"0A250B25", x"0C250D25", x"0E250F25",
		x"10251125", x"12251325", x"14251525", x"16251725", x"18251925", x"1A251B25", x"1C251D25", x"1E251F25",
		x"20252125", x"22252325", x"24252525", x"26252725", x"28252925", x"2A252B25", x"2C252D25", x"2E252F25",
		x"30253125", x"32253325", x"34253525", x"36253725", x"38253925", x"3A253B25", x"3C253D25", x"3E253F25",
		x"FFFFFFFF", x"FFFFFFFF", x"40254125", x"42254325", x"44254525", x"46254725", x"48254925", x"4A254B25",
		x"4C254D25", x"4E254F25", x"50255125", x"52255325", x"54255525", x"56255725", x"58255925", x"5A255B25",
		x"5C255D25", x"5E255F25", x"60256125", x"62256325", x"64256525", x"66256725", x"68256925", x"6A256B25",
		x"6C256D25", x"6E256F25", x"70257125", x"72257325", x"74257525", x"76257725", x"78257925", x"7A257B25",
		x"7C257D25", x"7E257F25", x"FFFFFFFF", x"FFFFFFFF", x"80258125", x"82258325", x"84258525", x"86258725",
		x"88258925", x"8A258B25", x"8C258D25", x"8E258F25", x"90259125", x"92259325", x"94259525", x"96259725",
		x"98259925", x"9A259B25", x"9C259D25", x"9E259F25", x"A025A125", x"A225A325", x"A425A525", x"A625A725",
		x"A825A925", x"AA25AB25", x"AC25AD25", x"AE25AF25", x"B025B125", x"B225B325", x"B425B525", x"B625B725",
		x"B825B925", x"BA25BB25", x"BC25BD25", x"BE25BF25", x"FFFFFFFF", x"FFFFFFFF", x"C025C125", x"C225C325",
		x"C425C525", x"C625C725", x"C825C925", x"CA25CB25", x"CC25CD25", x"CE25CF25", x"D025D125", x"D225D325",
		x"D425D525", x"D625D725", x"D825D925", x"DA25DB25", x"DC25DD25", x"DE25DF25", x"E025E125", x"E225E325",
		x"E425E525", x"E625E725", x"E825E925", x"EA25EB25", x"EC25ED25", x"EE25EF25", x"F025F125", x"F225F325",
		x"F425F525", x"F625F725", x"F825F925", x"FA25FB25", x"FC25FD25", x"FE25FF25", x"FFFFFFFF", x"FFFFFFFF",
		x"00260126", x"02260326", x"04260526", x"06260726", x"08260926", x"0A260B26", x"0C260D26", x"0E260F26",
		x"10261126", x"12261326", x"14261526", x"16261726", x"18261926", x"1A261B26", x"1C261D26", x"1E261F26",
		x"20262126", x"22262326", x"24262526", x"26262726", x"28262926", x"2A262B26", x"2C262D26", x"2E262F26",
		x"30263126", x"32263326", x"34263526", x"36263726", x"38263926", x"3A263B26", x"3C263D26", x"3E263F26",
		x"FFFFFFFF", x"FFFFFFFF", x"40264126", x"42264326", x"44264526", x"46264726", x"48264926", x"4A264B26",
		x"4C264D26", x"4E264F26", x"50265126", x"52265326", x"54265526", x"56265726", x"58265926", x"5A265B26",
		x"5C265D26", x"5E265F26", x"60266126", x"62266326", x"64266526", x"66266726", x"68266926", x"6A266B26",
		x"6C266D26", x"6E266F26", x"70267126", x"72267326", x"74267526", x"76267726", x"78267926", x"7A267B26",
		x"7C267D26", x"7E267F26", x"FFFFFFFF", x"FFFFFFFF", x"80268126", x"82268326", x"84268526", x"86268726",
		x"88268926", x"8A268B26", x"8C268D26", x"8E268F26", x"90269126", x"92269326", x"94269526", x"96269726",
		x"98269926", x"9A269B26", x"9C269D26", x"9E269F26", x"A026A126", x"A226A326", x"A426A526", x"A626A726",
		x"A826A926", x"AA26AB26", x"AC26AD26", x"AE26AF26", x"B026B126", x"B226B326", x"B426B526", x"B626B726",
		x"B826B926", x"BA26BB26", x"BC26BD26", x"BE26BF26", x"FFFFFFFF", x"FFFFFFFF", x"C026C126", x"C226C326",
		x"C426C526", x"C626C726", x"C826C926", x"CA26CB26", x"CC26CD26", x"CE26CF26", x"D026D126", x"D226D326",
		x"D426D526", x"D626D726", x"D826D926", x"DA26DB26", x"DC26DD26", x"DE26DF26", x"E026E126", x"E226E326",
		x"E426E526", x"E626E726", x"E826E926", x"EA26EB26", x"EC26ED26", x"EE26EF26", x"F026F126", x"F226F326",
		x"F426F526", x"F626F726", x"F826F926", x"FA26FB26", x"FC26FD26", x"FE26FF26", x"FFFFFFFF", x"FFFFFFFF",
		x"00270127", x"02270327", x"04270527", x"06270727", x"08270927", x"0A270B27", x"0C270D27", x"0E270F27",
		x"10271127", x"12271327", x"14271527", x"16271727", x"18271927", x"1A271B27", x"1C271D27", x"1E271F27",
		x"20272127", x"22272327", x"24272527", x"26272727", x"28272927", x"2A272B27", x"2C272D27", x"2E272F27",
		x"30273127", x"32273327", x"34273527", x"36273727", x"38273927", x"3A273B27", x"3C273D27", x"3E273F27",
		x"FFFFFFFF", x"FFFFFFFF", x"40274127", x"42274327", x"44274527", x"46274727", x"48274927", x"4A274B27",
		x"4C274D27", x"4E274F27", x"50275127", x"52275327", x"54275527", x"56275727", x"58275927", x"5A275B27",
		x"5C275D27", x"5E275F27", x"60276127", x"62276327", x"64276527", x"66276727", x"68276927", x"6A276B27",
		x"6C276D27", x"6E276F27", x"70277127", x"72277327", x"74277527", x"76277727", x"78277927", x"7A277B27",
		x"7C277D27", x"7E277F27", x"FFFFFFFF", x"FFFFFFFF", x"80278127", x"82278327", x"84278527", x"86278727",
		x"88278927", x"8A278B27", x"8C278D27", x"8E278F27", x"90279127", x"92279327", x"94279527", x"96279727",
		x"98279927", x"9A279B27", x"9C279D27", x"9E279F27", x"A027A127", x"A227A327", x"A427A527", x"A627A727",
		x"A827A927", x"AA27AB27", x"AC27AD27", x"AE27AF27", x"B027B127", x"B227B327", x"B427B527", x"B627B727",
		x"B827B927", x"BA27BB27", x"BC27BD27", x"BE27BF27", x"FFFFFFFF", x"FFFFFFFF", x"C027C127", x"C227C327",
		x"C427C527", x"C627C727", x"C827C927", x"CA27CB27", x"CC27CD27", x"CE27CF27", x"D027D127", x"D227D327",
		x"D427D527", x"D627D727", x"D827D927", x"DA27DB27", x"DC27DD27", x"DE27DF27", x"E027E127", x"E227E327",
		x"E427E527", x"E627E727", x"E827E927", x"EA27EB27", x"EC27ED27", x"EE27EF27", x"F027F127", x"F227F327",
		x"F427F527", x"F627F727", x"F827F927", x"FA27FB27", x"FC27FD27", x"FE27FF27", x"FFFFFFFF", x"FFFFFFFF",
		x"00280128", x"02280328", x"04280528", x"06280728", x"08280928", x"0A280B28", x"0C280D28", x"0E280F28",
		x"10281128", x"12281328", x"14281528", x"16281728", x"18281928", x"1A281B28", x"1C281D28", x"1E281F28",
		x"20282128", x"22282328", x"24282528", x"26282728", x"28282928", x"2A282B28", x"2C282D28", x"2E282F28",
		x"30283128", x"32283328", x"34283528", x"36283728", x"38283928", x"3A283B28", x"3C283D28", x"3E283F28",
		x"FFFFFFFF", x"FFFFFFFF", x"40284128", x"42284328", x"44284528", x"46284728", x"48284928", x"4A284B28",
		x"4C284D28", x"4E284F28", x"50285128", x"52285328", x"54285528", x"56285728", x"58285928", x"5A285B28",
		x"5C285D28", x"5E285F28", x"60286128", x"62286328", x"64286528", x"66286728", x"68286928", x"6A286B28",
		x"6C286D28", x"6E286F28", x"70287128", x"72287328", x"74287528", x"76287728", x"78287928", x"7A287B28",
		x"7C287D28", x"7E287F28", x"FFFFFFFF", x"FFFFFFFF", x"80288128", x"82288328", x"84288528", x"86288728",
		x"88288928", x"8A288B28", x"8C288D28", x"8E288F28", x"90289128", x"92289328", x"94289528", x"96289728",
		x"98289928", x"9A289B28", x"9C289D28", x"9E289F28", x"A028A128", x"A228A328", x"A428A528", x"A628A728",
		x"A828A928", x"AA28AB28", x"AC28AD28", x"AE28AF28", x"B028B128", x"B228B328", x"B428B528", x"B628B728",
		x"B828B928", x"BA28BB28", x"BC28BD28", x"BE28BF28", x"FFFFFFFF", x"FFFFFFFF", x"C028C128", x"C228C328",
		x"C428C528", x"C628C728", x"C828C928", x"CA28CB28", x"CC28CD28", x"CE28CF28", x"D028D128", x"D228D328",
		x"D428D528", x"D628D728", x"D828D928", x"DA28DB28", x"DC28DD28", x"DE28DF28", x"E028E128", x"E228E328",
		x"E428E528", x"E628E728", x"E828E928", x"EA28EB28", x"EC28ED28", x"EE28EF28", x"F028F128", x"F228F328",
		x"F428F528", x"F628F728", x"F828F928", x"FA28FB28", x"FC28FD28", x"FE28FF28", x"FFFFFFFF", x"FFFFFFFF",
		x"00290129", x"02290329", x"04290529", x"06290729", x"08290929", x"0A290B29", x"0C290D29", x"0E290F29",
		x"10291129", x"12291329", x"14291529", x"16291729", x"18291929", x"1A291B29", x"1C291D29", x"1E291F29",
		x"20292129", x"22292329", x"24292529", x"26292729", x"28292929", x"2A292B29", x"2C292D29", x"2E292F29",
		x"30293129", x"32293329", x"34293529", x"36293729", x"38293929", x"3A293B29", x"3C293D29", x"3E293F29",
		x"FFFFFFFF", x"FFFFFFFF", x"40294129", x"42294329", x"44294529", x"46294729", x"48294929", x"4A294B29",
		x"4C294D29", x"4E294F29", x"50295129", x"52295329", x"54295529", x"56295729", x"58295929", x"5A295B29",
		x"5C295D29", x"5E295F29", x"60296129", x"62296329", x"64296529", x"66296729", x"68296929", x"6A296B29",
		x"6C296D29", x"6E296F29", x"70297129", x"72297329", x"74297529", x"76297729", x"78297929", x"7A297B29",
		x"7C297D29", x"7E297F29", x"FFFFFFFF", x"FFFFFFFF", x"80298129", x"82298329", x"84298529", x"86298729",
		x"88298929", x"8A298B29", x"8C298D29", x"8E298F29", x"90299129", x"92299329", x"94299529", x"96299729",
		x"98299929", x"9A299B29", x"9C299D29", x"9E299F29", x"A029A129", x"A229A329", x"A429A529", x"A629A729",
		x"A829A929", x"AA29AB29", x"AC29AD29", x"AE29AF29", x"B029B129", x"B229B329", x"B429B529", x"B629B729",
		x"B829B929", x"BA29BB29", x"BC29BD29", x"BE29BF29", x"FFFFFFFF", x"FFFFFFFF", x"C029C129", x"C229C329",
		x"C429C529", x"C629C729", x"C829C929", x"CA29CB29", x"CC29CD29", x"CE29CF29", x"D029D129", x"D229D329",
		x"D429D529", x"D629D729", x"D829D929", x"DA29DB29", x"DC29DD29", x"DE29DF29", x"E029E129", x"E229E329",
		x"E429E529", x"E629E729", x"E829E929", x"EA29EB29", x"EC29ED29", x"EE29EF29", x"F029F129", x"F229F329",
		x"F429F529", x"F629F729", x"F829F929", x"FA29FB29", x"FC29FD29", x"FE29FF29", x"FFFFFFFF", x"FFFFFFFF",
		x"002A012A", x"022A032A", x"042A052A", x"062A072A", x"082A092A", x"0A2A0B2A", x"0C2A0D2A", x"0E2A0F2A",
		x"102A112A", x"122A132A", x"142A152A", x"162A172A", x"182A192A", x"1A2A1B2A", x"1C2A1D2A", x"1E2A1F2A",
		x"202A212A", x"222A232A", x"242A252A", x"262A272A", x"282A292A", x"2A2A2B2A", x"2C2A2D2A", x"2E2A2F2A",
		x"302A312A", x"322A332A", x"342A352A", x"362A372A", x"382A392A", x"3A2A3B2A", x"3C2A3D2A", x"3E2A3F2A",
		x"FFFFFFFF", x"FFFFFFFF", x"402A412A", x"422A432A", x"442A452A", x"462A472A", x"482A492A", x"4A2A4B2A",
		x"4C2A4D2A", x"4E2A4F2A", x"502A512A", x"522A532A", x"542A552A", x"562A572A", x"582A592A", x"5A2A5B2A",
		x"5C2A5D2A", x"5E2A5F2A", x"602A612A", x"622A632A", x"642A652A", x"662A672A", x"682A692A", x"6A2A6B2A",
		x"6C2A6D2A", x"6E2A6F2A", x"702A712A", x"722A732A", x"742A752A", x"762A772A", x"782A792A", x"7A2A7B2A",
		x"7C2A7D2A", x"7E2A7F2A", x"FFFFFFFF", x"FFFFFFFF", x"802A812A", x"822A832A", x"842A852A", x"862A872A",
		x"882A892A", x"8A2A8B2A", x"8C2A8D2A", x"8E2A8F2A", x"902A912A", x"922A932A", x"942A952A", x"962A972A",
		x"982A992A", x"9A2A9B2A", x"9C2A9D2A", x"9E2A9F2A", x"A02AA12A", x"A22AA32A", x"A42AA52A", x"A62AA72A",
		x"A82AA92A", x"AA2AAB2A", x"AC2AAD2A", x"AE2AAF2A", x"B02AB12A", x"B22AB32A", x"B42AB52A", x"B62AB72A",
		x"B82AB92A", x"BA2ABB2A", x"BC2ABD2A", x"BE2ABF2A", x"FFFFFFFF", x"FFFFFFFF", x"C02AC12A", x"C22AC32A",
		x"C42AC52A", x"C62AC72A", x"C82AC92A", x"CA2ACB2A", x"CC2ACD2A", x"CE2ACF2A", x"D02AD12A", x"D22AD32A",
		x"D42AD52A", x"D62AD72A", x"D82AD92A", x"DA2ADB2A", x"DC2ADD2A", x"DE2ADF2A", x"E02AE12A", x"E22AE32A",
		x"E42AE52A", x"E62AE72A", x"E82AE92A", x"EA2AEB2A", x"EC2AED2A", x"EE2AEF2A", x"F02AF12A", x"F22AF32A",
		x"F42AF52A", x"F62AF72A", x"F82AF92A", x"FA2AFB2A", x"FC2AFD2A", x"FE2AFF2A", x"FFFFFFFF", x"FFFFFFFF",
		x"002B012B", x"022B032B", x"042B052B", x"062B072B", x"082B092B", x"0A2B0B2B", x"0C2B0D2B", x"0E2B0F2B",
		x"102B112B", x"122B132B", x"142B152B", x"162B172B", x"182B192B", x"1A2B1B2B", x"1C2B1D2B", x"1E2B1F2B",
		x"202B212B", x"222B232B", x"242B252B", x"262B272B", x"282B292B", x"2A2B2B2B", x"2C2B2D2B", x"2E2B2F2B",
		x"302B312B", x"322B332B", x"342B352B", x"362B372B", x"382B392B", x"3A2B3B2B", x"3C2B3D2B", x"3E2B3F2B",
		x"FFFFFFFF", x"FFFFFFFF", x"402B412B", x"422B432B", x"442B452B", x"462B472B", x"482B492B", x"4A2B4B2B",
		x"4C2B4D2B", x"4E2B4F2B", x"502B512B", x"522B532B", x"542B552B", x"562B572B", x"582B592B", x"5A2B5B2B",
		x"5C2B5D2B", x"5E2B5F2B", x"602B612B", x"622B632B", x"642B652B", x"662B672B", x"682B692B", x"6A2B6B2B",
		x"6C2B6D2B", x"6E2B6F2B", x"702B712B", x"722B732B", x"742B752B", x"762B772B", x"782B792B", x"7A2B7B2B",
		x"7C2B7D2B", x"7E2B7F2B", x"FFFFFFFF", x"FFFFFFFF", x"802B812B", x"822B832B", x"842B852B", x"862B872B",
		x"882B892B", x"8A2B8B2B", x"8C2B8D2B", x"8E2B8F2B", x"902B912B", x"922B932B", x"942B952B", x"962B972B",
		x"982B992B", x"9A2B9B2B", x"9C2B9D2B", x"9E2B9F2B", x"A02BA12B", x"A22BA32B", x"A42BA52B", x"A62BA72B",
		x"A82BA92B", x"AA2BAB2B", x"AC2BAD2B", x"AE2BAF2B", x"B02BB12B", x"B22BB32B", x"B42BB52B", x"B62BB72B",
		x"B82BB92B", x"BA2BBB2B", x"BC2BBD2B", x"BE2BBF2B", x"FFFFFFFF", x"FFFFFFFF", x"C02BC12B", x"C22BC32B",
		x"C42BC52B", x"C62BC72B", x"C82BC92B", x"CA2BCB2B", x"CC2BCD2B", x"CE2BCF2B", x"D02BD12B", x"D22BD32B",
		x"D42BD52B", x"D62BD72B", x"D82BD92B", x"DA2BDB2B", x"DC2BDD2B", x"DE2BDF2B", x"E02BE12B", x"E22BE32B",
		x"E42BE52B", x"E62BE72B", x"E82BE92B", x"EA2BEB2B", x"EC2BED2B", x"EE2BEF2B", x"F02BF12B", x"F22BF32B",
		x"F42BF52B", x"F62BF72B", x"F82BF92B", x"FA2BFB2B", x"FC2BFD2B", x"FE2BFF2B", x"FFFFFFFF", x"FFFFFFFF",
		x"002C012C", x"022C032C", x"042C052C", x"062C072C", x"082C092C", x"0A2C0B2C", x"0C2C0D2C", x"0E2C0F2C",
		x"102C112C", x"122C132C", x"142C152C", x"162C172C", x"182C192C", x"1A2C1B2C", x"1C2C1D2C", x"1E2C1F2C",
		x"202C212C", x"222C232C", x"242C252C", x"262C272C", x"282C292C", x"2A2C2B2C", x"2C2C2D2C", x"2E2C2F2C",
		x"302C312C", x"322C332C", x"342C352C", x"362C372C", x"382C392C", x"3A2C3B2C", x"3C2C3D2C", x"3E2C3F2C",
		x"FFFFFFFF", x"FFFFFFFF", x"402C412C", x"422C432C", x"442C452C", x"462C472C", x"482C492C", x"4A2C4B2C",
		x"4C2C4D2C", x"4E2C4F2C", x"502C512C", x"522C532C", x"542C552C", x"562C572C", x"582C592C", x"5A2C5B2C",
		x"5C2C5D2C", x"5E2C5F2C", x"602C612C", x"622C632C", x"642C652C", x"662C672C", x"682C692C", x"6A2C6B2C",
		x"6C2C6D2C", x"6E2C6F2C", x"702C712C", x"722C732C", x"742C752C", x"762C772C", x"782C792C", x"7A2C7B2C",
		x"7C2C7D2C", x"7E2C7F2C", x"FFFFFFFF", x"FFFFFFFF", x"802C812C", x"822C832C", x"842C852C", x"862C872C",
		x"882C892C", x"8A2C8B2C", x"8C2C8D2C", x"8E2C8F2C", x"902C912C", x"922C932C", x"942C952C", x"962C972C",
		x"982C992C", x"9A2C9B2C", x"9C2C9D2C", x"9E2C9F2C", x"A02CA12C", x"A22CA32C", x"A42CA52C", x"A62CA72C",
		x"A82CA92C", x"AA2CAB2C", x"AC2CAD2C", x"AE2CAF2C", x"B02CB12C", x"B22CB32C", x"B42CB52C", x"B62CB72C",
		x"B82CB92C", x"BA2CBB2C", x"BC2CBD2C", x"BE2CBF2C", x"FFFFFFFF", x"FFFFFFFF", x"C02CC12C", x"C22CC32C",
		x"C42CC52C", x"C62CC72C", x"C82CC92C", x"CA2CCB2C", x"CC2CCD2C", x"CE2CCF2C", x"D02CD12C", x"D22CD32C",
		x"D42CD52C", x"D62CD72C", x"D82CD92C", x"DA2CDB2C", x"DC2CDD2C", x"DE2CDF2C", x"E02CE12C", x"E22CE32C",
		x"E42CE52C", x"E62CE72C", x"E82CE92C", x"EA2CEB2C", x"EC2CED2C", x"EE2CEF2C", x"F02CF12C", x"F22CF32C",
		x"F42CF52C", x"F62CF72C", x"F82CF92C", x"FA2CFB2C", x"FC2CFD2C", x"FE2CFF2C", x"FFFFFFFF", x"FFFFFFFF",
		x"002D012D", x"022D032D", x"042D052D", x"062D072D", x"082D092D", x"0A2D0B2D", x"0C2D0D2D", x"0E2D0F2D",
		x"102D112D", x"122D132D", x"142D152D", x"162D172D", x"182D192D", x"1A2D1B2D", x"1C2D1D2D", x"1E2D1F2D",
		x"202D212D", x"222D232D", x"242D252D", x"262D272D", x"282D292D", x"2A2D2B2D", x"2C2D2D2D", x"2E2D2F2D",
		x"302D312D", x"322D332D", x"342D352D", x"362D372D", x"382D392D", x"3A2D3B2D", x"3C2D3D2D", x"3E2D3F2D",
		x"FFFFFFFF", x"FFFFFFFF", x"402D412D", x"422D432D", x"442D452D", x"462D472D", x"482D492D", x"4A2D4B2D",
		x"4C2D4D2D", x"4E2D4F2D", x"502D512D", x"522D532D", x"542D552D", x"562D572D", x"582D592D", x"5A2D5B2D",
		x"5C2D5D2D", x"5E2D5F2D", x"602D612D", x"622D632D", x"642D652D", x"662D672D", x"682D692D", x"6A2D6B2D",
		x"6C2D6D2D", x"6E2D6F2D", x"702D712D", x"722D732D", x"742D752D", x"762D772D", x"782D792D", x"7A2D7B2D",
		x"7C2D7D2D", x"7E2D7F2D", x"FFFFFFFF", x"FFFFFFFF", x"802D812D", x"822D832D", x"842D852D", x"862D872D",
		x"882D892D", x"8A2D8B2D", x"8C2D8D2D", x"8E2D8F2D", x"902D912D", x"922D932D", x"942D952D", x"962D972D",
		x"982D992D", x"9A2D9B2D", x"9C2D9D2D", x"9E2D9F2D", x"A02DA12D", x"A22DA32D", x"A42DA52D", x"A62DA72D",
		x"A82DA92D", x"AA2DAB2D", x"AC2DAD2D", x"AE2DAF2D", x"B02DB12D", x"B22DB32D", x"B42DB52D", x"B62DB72D",
		x"B82DB92D", x"BA2DBB2D", x"BC2DBD2D", x"BE2DBF2D", x"FFFFFFFF", x"FFFFFFFF", x"C02DC12D", x"C22DC32D",
		x"C42DC52D", x"C62DC72D", x"C82DC92D", x"CA2DCB2D", x"CC2DCD2D", x"CE2DCF2D", x"D02DD12D", x"D22DD32D",
		x"D42DD52D", x"D62DD72D", x"D82DD92D", x"DA2DDB2D", x"DC2DDD2D", x"DE2DDF2D", x"E02DE12D", x"E22DE32D",
		x"E42DE52D", x"E62DE72D", x"E82DE92D", x"EA2DEB2D", x"EC2DED2D", x"EE2DEF2D", x"F02DF12D", x"F22DF32D",
		x"F42DF52D", x"F62DF72D", x"F82DF92D", x"FA2DFB2D", x"FC2DFD2D", x"FE2DFF2D", x"FFFFFFFF", x"FFFFFFFF",
		x"002E012E", x"022E032E", x"042E052E", x"062E072E", x"082E092E", x"0A2E0B2E", x"0C2E0D2E", x"0E2E0F2E",
		x"102E112E", x"122E132E", x"142E152E", x"162E172E", x"182E192E", x"1A2E1B2E", x"1C2E1D2E", x"1E2E1F2E",
		x"202E212E", x"222E232E", x"242E252E", x"262E272E", x"282E292E", x"2A2E2B2E", x"2C2E2D2E", x"2E2E2F2E",
		x"302E312E", x"322E332E", x"342E352E", x"362E372E", x"382E392E", x"3A2E3B2E", x"3C2E3D2E", x"3E2E3F2E",
		x"FFFFFFFF", x"FFFFFFFF", x"402E412E", x"422E432E", x"442E452E", x"462E472E", x"482E492E", x"4A2E4B2E",
		x"4C2E4D2E", x"4E2E4F2E", x"502E512E", x"522E532E", x"542E552E", x"562E572E", x"582E592E", x"5A2E5B2E",
		x"5C2E5D2E", x"5E2E5F2E", x"602E612E", x"622E632E", x"642E652E", x"662E672E", x"682E692E", x"6A2E6B2E",
		x"6C2E6D2E", x"6E2E6F2E", x"702E712E", x"722E732E", x"742E752E", x"762E772E", x"782E792E", x"7A2E7B2E",
		x"7C2E7D2E", x"7E2E7F2E", x"FFFFFFFF", x"FFFFFFFF", x"802E812E", x"822E832E", x"842E852E", x"862E872E",
		x"882E892E", x"8A2E8B2E", x"8C2E8D2E", x"8E2E8F2E", x"902E912E", x"922E932E", x"942E952E", x"962E972E",
		x"982E992E", x"9A2E9B2E", x"9C2E9D2E", x"9E2E9F2E", x"A02EA12E", x"A22EA32E", x"A42EA52E", x"A62EA72E",
		x"A82EA92E", x"AA2EAB2E", x"AC2EAD2E", x"AE2EAF2E", x"B02EB12E", x"B22EB32E", x"B42EB52E", x"B62EB72E",
		x"B82EB92E", x"BA2EBB2E", x"BC2EBD2E", x"BE2EBF2E", x"FFFFFFFF", x"FFFFFFFF", x"C02EC12E", x"C22EC32E",
		x"C42EC52E", x"C62EC72E", x"C82EC92E", x"CA2ECB2E", x"CC2ECD2E", x"CE2ECF2E", x"D02ED12E", x"D22ED32E",
		x"D42ED52E", x"D62ED72E", x"D82ED92E", x"DA2EDB2E", x"DC2EDD2E", x"DE2EDF2E", x"E02EE12E", x"E22EE32E",
		x"E42EE52E", x"E62EE72E", x"E82EE92E", x"EA2EEB2E", x"EC2EED2E", x"EE2EEF2E", x"F02EF12E", x"F22EF32E",
		x"F42EF52E", x"F62EF72E", x"F82EF92E", x"FA2EFB2E", x"FC2EFD2E", x"FE2EFF2E", x"FFFFFFFF", x"FFFFFFFF",
		x"002F012F", x"022F032F", x"042F052F", x"062F072F", x"082F092F", x"0A2F0B2F", x"0C2F0D2F", x"0E2F0F2F",
		x"102F112F", x"122F132F", x"142F152F", x"162F172F", x"182F192F", x"1A2F1B2F", x"1C2F1D2F", x"1E2F1F2F",
		x"202F212F", x"222F232F", x"242F252F", x"262F272F", x"282F292F", x"2A2F2B2F", x"2C2F2D2F", x"2E2F2F2F",
		x"302F312F", x"322F332F", x"342F352F", x"362F372F", x"382F392F", x"3A2F3B2F", x"3C2F3D2F", x"3E2F3F2F",
		x"FFFFFFFF", x"FFFFFFFF", x"402F412F", x"422F432F", x"442F452F", x"462F472F", x"482F492F", x"4A2F4B2F",
		x"4C2F4D2F", x"4E2F4F2F", x"502F512F", x"522F532F", x"542F552F", x"562F572F", x"582F592F", x"5A2F5B2F",
		x"5C2F5D2F", x"5E2F5F2F", x"602F612F", x"622F632F", x"642F652F", x"662F672F", x"682F692F", x"6A2F6B2F",
		x"6C2F6D2F", x"6E2F6F2F", x"702F712F", x"722F732F", x"742F752F", x"762F772F", x"782F792F", x"7A2F7B2F",
		x"7C2F7D2F", x"7E2F7F2F", x"FFFFFFFF", x"FFFFFFFF", x"802F812F", x"822F832F", x"842F852F", x"862F872F",
		x"882F892F", x"8A2F8B2F", x"8C2F8D2F", x"8E2F8F2F", x"902F912F", x"922F932F", x"942F952F", x"962F972F",
		x"982F992F", x"9A2F9B2F", x"9C2F9D2F", x"9E2F9F2F", x"A02FA12F", x"A22FA32F", x"A42FA52F", x"A62FA72F",
		x"A82FA92F", x"AA2FAB2F", x"AC2FAD2F", x"AE2FAF2F", x"B02FB12F", x"B22FB32F", x"B42FB52F", x"B62FB72F",
		x"B82FB92F", x"BA2FBB2F", x"BC2FBD2F", x"BE2FBF2F", x"FFFFFFFF", x"FFFFFFFF", x"C02FC12F", x"C22FC32F",
		x"C42FC52F", x"C62FC72F", x"C82FC92F", x"CA2FCB2F", x"CC2FCD2F", x"CE2FCF2F", x"D02FD12F", x"D22FD32F",
		x"D42FD52F", x"D62FD72F", x"D82FD92F", x"DA2FDB2F", x"DC2FDD2F", x"DE2FDF2F", x"E02FE12F", x"E22FE32F",
		x"E42FE52F", x"E62FE72F", x"E82FE92F", x"EA2FEB2F", x"EC2FED2F", x"EE2FEF2F", x"F02FF12F", x"F22FF32F",
		x"F42FF52F", x"F62FF72F", x"F82FF92F", x"FA2FFB2F", x"FC2FFD2F", x"FE2FFF2F", x"FFFFFFFF", x"FFFFFFFF",
		x"00300130", x"02300330", x"04300530", x"06300730", x"08300930", x"0A300B30", x"0C300D30", x"0E300F30",
		x"10301130", x"12301330", x"14301530", x"16301730", x"18301930", x"1A301B30", x"1C301D30", x"1E301F30",
		x"20302130", x"22302330", x"24302530", x"26302730", x"28302930", x"2A302B30", x"2C302D30", x"2E302F30",
		x"30303130", x"32303330", x"34303530", x"36303730", x"38303930", x"3A303B30", x"3C303D30", x"3E303F30",
		x"FFFFFFFF", x"FFFFFFFF", x"40304130", x"42304330", x"44304530", x"46304730", x"48304930", x"4A304B30",
		x"4C304D30", x"4E304F30", x"50305130", x"52305330", x"54305530", x"56305730", x"58305930", x"5A305B30",
		x"5C305D30", x"5E305F30", x"60306130", x"62306330", x"64306530", x"66306730", x"68306930", x"6A306B30",
		x"6C306D30", x"6E306F30", x"70307130", x"72307330", x"74307530", x"76307730", x"78307930", x"7A307B30",
		x"7C307D30", x"7E307F30", x"FFFFFFFF", x"FFFFFFFF", x"80308130", x"82308330", x"84308530", x"86308730",
		x"88308930", x"8A308B30", x"8C308D30", x"8E308F30", x"90309130", x"92309330", x"94309530", x"96309730",
		x"98309930", x"9A309B30", x"9C309D30", x"9E309F30", x"A030A130", x"A230A330", x"A430A530", x"A630A730",
		x"A830A930", x"AA30AB30", x"AC30AD30", x"AE30AF30", x"B030B130", x"B230B330", x"B430B530", x"B630B730",
		x"B830B930", x"BA30BB30", x"BC30BD30", x"BE30BF30", x"FFFFFFFF", x"FFFFFFFF", x"C030C130", x"C230C330",
		x"C430C530", x"C630C730", x"C830C930", x"CA30CB30", x"CC30CD30", x"CE30CF30", x"D030D130", x"D230D330",
		x"D430D530", x"D630D730", x"D830D930", x"DA30DB30", x"DC30DD30", x"DE30DF30", x"E030E130", x"E230E330",
		x"E430E530", x"E630E730", x"E830E930", x"EA30EB30", x"EC30ED30", x"EE30EF30", x"F030F130", x"F230F330",
		x"F430F530", x"F630F730", x"F830F930", x"FA30FB30", x"FC30FD30", x"FE30FF30", x"FFFFFFFF", x"FFFFFFFF",
		x"00310131", x"02310331", x"04310531", x"06310731", x"08310931", x"0A310B31", x"0C310D31", x"0E310F31",
		x"10311131", x"12311331", x"14311531", x"16311731", x"18311931", x"1A311B31", x"1C311D31", x"1E311F31",
		x"20312131", x"22312331", x"24312531", x"26312731", x"28312931", x"2A312B31", x"2C312D31", x"2E312F31",
		x"30313131", x"32313331", x"34313531", x"36313731", x"38313931", x"3A313B31", x"3C313D31", x"3E313F31",
		x"FFFFFFFF", x"FFFFFFFF", x"40314131", x"42314331", x"44314531", x"46314731", x"48314931", x"4A314B31",
		x"4C314D31", x"4E314F31", x"50315131", x"52315331", x"54315531", x"56315731", x"58315931", x"5A315B31",
		x"5C315D31", x"5E315F31", x"60316131", x"62316331", x"64316531", x"66316731", x"68316931", x"6A316B31",
		x"6C316D31", x"6E316F31", x"70317131", x"72317331", x"74317531", x"76317731", x"78317931", x"7A317B31",
		x"7C317D31", x"7E317F31", x"FFFFFFFF", x"FFFFFFFF", x"80318131", x"82318331", x"84318531", x"86318731",
		x"88318931", x"8A318B31", x"8C318D31", x"8E318F31", x"90319131", x"92319331", x"94319531", x"96319731",
		x"98319931", x"9A319B31", x"9C319D31", x"9E319F31", x"A031A131", x"A231A331", x"A431A531", x"A631A731",
		x"A831A931", x"AA31AB31", x"AC31AD31", x"AE31AF31", x"B031B131", x"B231B331", x"B431B531", x"B631B731",
		x"B831B931", x"BA31BB31", x"BC31BD31", x"BE31BF31", x"FFFFFFFF", x"FFFFFFFF", x"C031C131", x"C231C331",
		x"C431C531", x"C631C731", x"C831C931", x"CA31CB31", x"CC31CD31", x"CE31CF31", x"D031D131", x"D231D331",
		x"D431D531", x"D631D731", x"D831D931", x"DA31DB31", x"DC31DD31", x"DE31DF31", x"E031E131", x"E231E331",
		x"E431E531", x"E631E731", x"E831E931", x"EA31EB31", x"EC31ED31", x"EE31EF31", x"F031F131", x"F231F331",
		x"F431F531", x"F631F731", x"F831F931", x"FA31FB31", x"FC31FD31", x"FE31FF31", x"FFFFFFFF", x"FFFFFFFF",
		x"00320132", x"02320332", x"04320532", x"06320732", x"08320932", x"0A320B32", x"0C320D32", x"0E320F32",
		x"10321132", x"12321332", x"14321532", x"16321732", x"18321932", x"1A321B32", x"1C321D32", x"1E321F32",
		x"20322132", x"22322332", x"24322532", x"26322732", x"28322932", x"2A322B32", x"2C322D32", x"2E322F32",
		x"30323132", x"32323332", x"34323532", x"36323732", x"38323932", x"3A323B32", x"3C323D32", x"3E323F32",
		x"FFFFFFFF", x"FFFFFFFF", x"40324132", x"42324332", x"44324532", x"46324732", x"48324932", x"4A324B32",
		x"4C324D32", x"4E324F32", x"50325132", x"52325332", x"54325532", x"56325732", x"58325932", x"5A325B32",
		x"5C325D32", x"5E325F32", x"60326132", x"62326332", x"64326532", x"66326732", x"68326932", x"6A326B32",
		x"6C326D32", x"6E326F32", x"70327132", x"72327332", x"74327532", x"76327732", x"78327932", x"7A327B32",
		x"7C327D32", x"7E327F32", x"FFFFFFFF", x"FFFFFFFF", x"80328132", x"82328332", x"84328532", x"86328732",
		x"88328932", x"8A328B32", x"8C328D32", x"8E328F32", x"90329132", x"92329332", x"94329532", x"96329732",
		x"98329932", x"9A329B32", x"9C329D32", x"9E329F32", x"A032A132", x"A232A332", x"A432A532", x"A632A732",
		x"A832A932", x"AA32AB32", x"AC32AD32", x"AE32AF32", x"B032B132", x"B232B332", x"B432B532", x"B632B732",
		x"B832B932", x"BA32BB32", x"BC32BD32", x"BE32BF32", x"FFFFFFFF", x"FFFFFFFF", x"C032C132", x"C232C332",
		x"C432C532", x"C632C732", x"C832C932", x"CA32CB32", x"CC32CD32", x"CE32CF32", x"D032D132", x"D232D332",
		x"D432D532", x"D632D732", x"D832D932", x"DA32DB32", x"DC32DD32", x"DE32DF32", x"E032E132", x"E232E332",
		x"E432E532", x"E632E732", x"E832E932", x"EA32EB32", x"EC32ED32", x"EE32EF32", x"F032F132", x"F232F332",
		x"F432F532", x"F632F732", x"F832F932", x"FA32FB32", x"FC32FD32", x"FE32FF32", x"FFFFFFFF", x"FFFFFFFF",
		x"00330133", x"02330333", x"04330533", x"06330733", x"08330933", x"0A330B33", x"0C330D33", x"0E330F33",
		x"10331133", x"12331333", x"14331533", x"16331733", x"18331933", x"1A331B33", x"1C331D33", x"1E331F33",
		x"20332133", x"22332333", x"24332533", x"26332733", x"28332933", x"2A332B33", x"2C332D33", x"2E332F33",
		x"30333133", x"32333333", x"34333533", x"36333733", x"38333933", x"3A333B33", x"3C333D33", x"3E333F33",
		x"FFFFFFFF", x"FFFFFFFF", x"40334133", x"42334333", x"44334533", x"46334733", x"48334933", x"4A334B33",
		x"4C334D33", x"4E334F33", x"50335133", x"52335333", x"54335533", x"56335733", x"58335933", x"5A335B33",
		x"5C335D33", x"5E335F33", x"60336133", x"62336333", x"64336533", x"66336733", x"68336933", x"6A336B33",
		x"6C336D33", x"6E336F33", x"70337133", x"72337333", x"74337533", x"76337733", x"78337933", x"7A337B33",
		x"7C337D33", x"7E337F33", x"FFFFFFFF", x"FFFFFFFF", x"80338133", x"82338333", x"84338533", x"86338733",
		x"88338933", x"8A338B33", x"8C338D33", x"8E338F33", x"90339133", x"92339333", x"94339533", x"96339733",
		x"98339933", x"9A339B33", x"9C339D33", x"9E339F33", x"A033A133", x"A233A333", x"A433A533", x"A633A733",
		x"A833A933", x"AA33AB33", x"AC33AD33", x"AE33AF33", x"B033B133", x"B233B333", x"B433B533", x"B633B733",
		x"B833B933", x"BA33BB33", x"BC33BD33", x"BE33BF33", x"FFFFFFFF", x"FFFFFFFF", x"C033C133", x"C233C333",
		x"C433C533", x"C633C733", x"C833C933", x"CA33CB33", x"CC33CD33", x"CE33CF33", x"D033D133", x"D233D333",
		x"D433D533", x"D633D733", x"D833D933", x"DA33DB33", x"DC33DD33", x"DE33DF33", x"E033E133", x"E233E333",
		x"E433E533", x"E633E733", x"E833E933", x"EA33EB33", x"EC33ED33", x"EE33EF33", x"F033F133", x"F233F333",
		x"F433F533", x"F633F733", x"F833F933", x"FA33FB33", x"FC33FD33", x"FE33FF33", x"FFFFFFFF", x"FFFFFFFF",
		x"00340134", x"02340334", x"04340534", x"06340734", x"08340934", x"0A340B34", x"0C340D34", x"0E340F34",
		x"10341134", x"12341334", x"14341534", x"16341734", x"18341934", x"1A341B34", x"1C341D34", x"1E341F34",
		x"20342134", x"22342334", x"24342534", x"26342734", x"28342934", x"2A342B34", x"2C342D34", x"2E342F34",
		x"30343134", x"32343334", x"34343534", x"36343734", x"38343934", x"3A343B34", x"3C343D34", x"3E343F34",
		x"FFFFFFFF", x"FFFFFFFF", x"40344134", x"42344334", x"44344534", x"46344734", x"48344934", x"4A344B34",
		x"4C344D34", x"4E344F34", x"50345134", x"52345334", x"54345534", x"56345734", x"58345934", x"5A345B34",
		x"5C345D34", x"5E345F34", x"60346134", x"62346334", x"64346534", x"66346734", x"68346934", x"6A346B34",
		x"6C346D34", x"6E346F34", x"70347134", x"72347334", x"74347534", x"76347734", x"78347934", x"7A347B34",
		x"7C347D34", x"7E347F34", x"FFFFFFFF", x"FFFFFFFF", x"80348134", x"82348334", x"84348534", x"86348734",
		x"88348934", x"8A348B34", x"8C348D34", x"8E348F34", x"90349134", x"92349334", x"94349534", x"96349734",
		x"98349934", x"9A349B34", x"9C349D34", x"9E349F34", x"A034A134", x"A234A334", x"A434A534", x"A634A734",
		x"A834A934", x"AA34AB34", x"AC34AD34", x"AE34AF34", x"B034B134", x"B234B334", x"B434B534", x"B634B734",
		x"B834B934", x"BA34BB34", x"BC34BD34", x"BE34BF34", x"FFFFFFFF", x"FFFFFFFF", x"C034C134", x"C234C334",
		x"C434C534", x"C634C734", x"C834C934", x"CA34CB34", x"CC34CD34", x"CE34CF34", x"D034D134", x"D234D334",
		x"D434D534", x"D634D734", x"D834D934", x"DA34DB34", x"DC34DD34", x"DE34DF34", x"E034E134", x"E234E334",
		x"E434E534", x"E634E734", x"E834E934", x"EA34EB34", x"EC34ED34", x"EE34EF34", x"F034F134", x"F234F334",
		x"F434F534", x"F634F734", x"F834F934", x"FA34FB34", x"FC34FD34", x"FE34FF34", x"FFFFFFFF", x"FFFFFFFF",
		x"00350135", x"02350335", x"04350535", x"06350735", x"08350935", x"0A350B35", x"0C350D35", x"0E350F35",
		x"10351135", x"12351335", x"14351535", x"16351735", x"18351935", x"1A351B35", x"1C351D35", x"1E351F35",
		x"20352135", x"22352335", x"24352535", x"26352735", x"28352935", x"2A352B35", x"2C352D35", x"2E352F35",
		x"30353135", x"32353335", x"34353535", x"36353735", x"38353935", x"3A353B35", x"3C353D35", x"3E353F35",
		x"FFFFFFFF", x"FFFFFFFF", x"40354135", x"42354335", x"44354535", x"46354735", x"48354935", x"4A354B35",
		x"4C354D35", x"4E354F35", x"50355135", x"52355335", x"54355535", x"56355735", x"58355935", x"5A355B35",
		x"5C355D35", x"5E355F35", x"60356135", x"62356335", x"64356535", x"66356735", x"68356935", x"6A356B35",
		x"6C356D35", x"6E356F35", x"70357135", x"72357335", x"74357535", x"76357735", x"78357935", x"7A357B35",
		x"7C357D35", x"7E357F35", x"FFFFFFFF", x"FFFFFFFF", x"80358135", x"82358335", x"84358535", x"86358735",
		x"88358935", x"8A358B35", x"8C358D35", x"8E358F35", x"90359135", x"92359335", x"94359535", x"96359735",
		x"98359935", x"9A359B35", x"9C359D35", x"9E359F35", x"A035A135", x"A235A335", x"A435A535", x"A635A735",
		x"A835A935", x"AA35AB35", x"AC35AD35", x"AE35AF35", x"B035B135", x"B235B335", x"B435B535", x"B635B735",
		x"B835B935", x"BA35BB35", x"BC35BD35", x"BE35BF35", x"FFFFFFFF", x"FFFFFFFF", x"C035C135", x"C235C335",
		x"C435C535", x"C635C735", x"C835C935", x"CA35CB35", x"CC35CD35", x"CE35CF35", x"D035D135", x"D235D335",
		x"D435D535", x"D635D735", x"D835D935", x"DA35DB35", x"DC35DD35", x"DE35DF35", x"E035E135", x"E235E335",
		x"E435E535", x"E635E735", x"E835E935", x"EA35EB35", x"EC35ED35", x"EE35EF35", x"F035F135", x"F235F335",
		x"F435F535", x"F635F735", x"F835F935", x"FA35FB35", x"FC35FD35", x"FE35FF35", x"FFFFFFFF", x"FFFFFFFF",
		x"00360136", x"02360336", x"04360536", x"06360736", x"08360936", x"0A360B36", x"0C360D36", x"0E360F36",
		x"10361136", x"12361336", x"14361536", x"16361736", x"18361936", x"1A361B36", x"1C361D36", x"1E361F36",
		x"20362136", x"22362336", x"24362536", x"26362736", x"28362936", x"2A362B36", x"2C362D36", x"2E362F36",
		x"30363136", x"32363336", x"34363536", x"36363736", x"38363936", x"3A363B36", x"3C363D36", x"3E363F36",
		x"FFFFFFFF", x"FFFFFFFF", x"40364136", x"42364336", x"44364536", x"46364736", x"48364936", x"4A364B36",
		x"4C364D36", x"4E364F36", x"50365136", x"52365336", x"54365536", x"56365736", x"58365936", x"5A365B36",
		x"5C365D36", x"5E365F36", x"60366136", x"62366336", x"64366536", x"66366736", x"68366936", x"6A366B36",
		x"6C366D36", x"6E366F36", x"70367136", x"72367336", x"74367536", x"76367736", x"78367936", x"7A367B36",
		x"7C367D36", x"7E367F36", x"FFFFFFFF", x"FFFFFFFF", x"80368136", x"82368336", x"84368536", x"86368736",
		x"88368936", x"8A368B36", x"8C368D36", x"8E368F36", x"90369136", x"92369336", x"94369536", x"96369736",
		x"98369936", x"9A369B36", x"9C369D36", x"9E369F36", x"A036A136", x"A236A336", x"A436A536", x"A636A736",
		x"A836A936", x"AA36AB36", x"AC36AD36", x"AE36AF36", x"B036B136", x"B236B336", x"B436B536", x"B636B736",
		x"B836B936", x"BA36BB36", x"BC36BD36", x"BE36BF36", x"FFFFFFFF", x"FFFFFFFF", x"C036C136", x"C236C336",
		x"C436C536", x"C636C736", x"C836C936", x"CA36CB36", x"CC36CD36", x"CE36CF36", x"D036D136", x"D236D336",
		x"D436D536", x"D636D736", x"D836D936", x"DA36DB36", x"DC36DD36", x"DE36DF36", x"E036E136", x"E236E336",
		x"E436E536", x"E636E736", x"E836E936", x"EA36EB36", x"EC36ED36", x"EE36EF36", x"F036F136", x"F236F336",
		x"F436F536", x"F636F736", x"F836F936", x"FA36FB36", x"FC36FD36", x"FE36FF36", x"FFFFFFFF", x"FFFFFFFF",
		x"00370137", x"02370337", x"04370537", x"06370737", x"08370937", x"0A370B37", x"0C370D37", x"0E370F37",
		x"10371137", x"12371337", x"14371537", x"16371737", x"18371937", x"1A371B37", x"1C371D37", x"1E371F37",
		x"20372137", x"22372337", x"24372537", x"26372737", x"28372937", x"2A372B37", x"2C372D37", x"2E372F37",
		x"30373137", x"32373337", x"34373537", x"36373737", x"38373937", x"3A373B37", x"3C373D37", x"3E373F37",
		x"FFFFFFFF", x"FFFFFFFF", x"40374137", x"42374337", x"44374537", x"46374737", x"48374937", x"4A374B37",
		x"4C374D37", x"4E374F37", x"50375137", x"52375337", x"54375537", x"56375737", x"58375937", x"5A375B37",
		x"5C375D37", x"5E375F37", x"60376137", x"62376337", x"64376537", x"66376737", x"68376937", x"6A376B37",
		x"6C376D37", x"6E376F37", x"70377137", x"72377337", x"74377537", x"76377737", x"78377937", x"7A377B37",
		x"7C377D37", x"7E377F37", x"FFFFFFFF", x"FFFFFFFF", x"80378137", x"82378337", x"84378537", x"86378737",
		x"88378937", x"8A378B37", x"8C378D37", x"8E378F37", x"90379137", x"92379337", x"94379537", x"96379737",
		x"98379937", x"9A379B37", x"9C379D37", x"9E379F37", x"A037A137", x"A237A337", x"A437A537", x"A637A737",
		x"A837A937", x"AA37AB37", x"AC37AD37", x"AE37AF37", x"B037B137", x"B237B337", x"B437B537", x"B637B737",
		x"B837B937", x"BA37BB37", x"BC37BD37", x"BE37BF37", x"FFFFFFFF", x"FFFFFFFF", x"C037C137", x"C237C337",
		x"C437C537", x"C637C737", x"C837C937", x"CA37CB37", x"CC37CD37", x"CE37CF37", x"D037D137", x"D237D337",
		x"D437D537", x"D637D737", x"D837D937", x"DA37DB37", x"DC37DD37", x"DE37DF37", x"E037E137", x"E237E337",
		x"E437E537", x"E637E737", x"E837E937", x"EA37EB37", x"EC37ED37", x"EE37EF37", x"F037F137", x"F237F337",
		x"F437F537", x"F637F737", x"F837F937", x"FA37FB37", x"FC37FD37", x"FE37FF37", x"FFFFFFFF", x"FFFFFFFF",
		x"00380138", x"02380338", x"04380538", x"06380738", x"08380938", x"0A380B38", x"0C380D38", x"0E380F38",
		x"10381138", x"12381338", x"14381538", x"16381738", x"18381938", x"1A381B38", x"1C381D38", x"1E381F38",
		x"20382138", x"22382338", x"24382538", x"26382738", x"28382938", x"2A382B38", x"2C382D38", x"2E382F38",
		x"30383138", x"32383338", x"34383538", x"36383738", x"38383938", x"3A383B38", x"3C383D38", x"3E383F38",
		x"FFFFFFFF", x"FFFFFFFF", x"40384138", x"42384338", x"44384538", x"46384738", x"48384938", x"4A384B38",
		x"4C384D38", x"4E384F38", x"50385138", x"52385338", x"54385538", x"56385738", x"58385938", x"5A385B38",
		x"5C385D38", x"5E385F38", x"60386138", x"62386338", x"64386538", x"66386738", x"68386938", x"6A386B38",
		x"6C386D38", x"6E386F38", x"70387138", x"72387338", x"74387538", x"76387738", x"78387938", x"7A387B38",
		x"7C387D38", x"7E387F38", x"FFFFFFFF", x"FFFFFFFF", x"80388138", x"82388338", x"84388538", x"86388738",
		x"88388938", x"8A388B38", x"8C388D38", x"8E388F38", x"90389138", x"92389338", x"94389538", x"96389738",
		x"98389938", x"9A389B38", x"9C389D38", x"9E389F38", x"A038A138", x"A238A338", x"A438A538", x"A638A738",
		x"A838A938", x"AA38AB38", x"AC38AD38", x"AE38AF38", x"B038B138", x"B238B338", x"B438B538", x"B638B738",
		x"B838B938", x"BA38BB38", x"BC38BD38", x"BE38BF38", x"FFFFFFFF", x"FFFFFFFF", x"C038C138", x"C238C338",
		x"C438C538", x"C638C738", x"C838C938", x"CA38CB38", x"CC38CD38", x"CE38CF38", x"D038D138", x"D238D338",
		x"D438D538", x"D638D738", x"D838D938", x"DA38DB38", x"DC38DD38", x"DE38DF38", x"E038E138", x"E238E338",
		x"E438E538", x"E638E738", x"E838E938", x"EA38EB38", x"EC38ED38", x"EE38EF38", x"F038F138", x"F238F338",
		x"F438F538", x"F638F738", x"F838F938", x"FA38FB38", x"FC38FD38", x"FE38FF38", x"FFFFFFFF", x"FFFFFFFF",
		x"00390139", x"02390339", x"04390539", x"06390739", x"08390939", x"0A390B39", x"0C390D39", x"0E390F39",
		x"10391139", x"12391339", x"14391539", x"16391739", x"18391939", x"1A391B39", x"1C391D39", x"1E391F39",
		x"20392139", x"22392339", x"24392539", x"26392739", x"28392939", x"2A392B39", x"2C392D39", x"2E392F39",
		x"30393139", x"32393339", x"34393539", x"36393739", x"38393939", x"3A393B39", x"3C393D39", x"3E393F39",
		x"FFFFFFFF", x"FFFFFFFF", x"40394139", x"42394339", x"44394539", x"46394739", x"48394939", x"4A394B39",
		x"4C394D39", x"4E394F39", x"50395139", x"52395339", x"54395539", x"56395739", x"58395939", x"5A395B39",
		x"5C395D39", x"5E395F39", x"60396139", x"62396339", x"64396539", x"66396739", x"68396939", x"6A396B39",
		x"6C396D39", x"6E396F39", x"70397139", x"72397339", x"74397539", x"76397739", x"78397939", x"7A397B39",
		x"7C397D39", x"7E397F39", x"FFFFFFFF", x"FFFFFFFF", x"80398139", x"82398339", x"84398539", x"86398739",
		x"88398939", x"8A398B39", x"8C398D39", x"8E398F39", x"90399139", x"92399339", x"94399539", x"96399739",
		x"98399939", x"9A399B39", x"9C399D39", x"9E399F39", x"A039A139", x"A239A339", x"A439A539", x"A639A739",
		x"A839A939", x"AA39AB39", x"AC39AD39", x"AE39AF39", x"B039B139", x"B239B339", x"B439B539", x"B639B739",
		x"B839B939", x"BA39BB39", x"BC39BD39", x"BE39BF39", x"FFFFFFFF", x"FFFFFFFF", x"C039C139", x"C239C339",
		x"C439C539", x"C639C739", x"C839C939", x"CA39CB39", x"CC39CD39", x"CE39CF39", x"D039D139", x"D239D339",
		x"D439D539", x"D639D739", x"D839D939", x"DA39DB39", x"DC39DD39", x"DE39DF39", x"E039E139", x"E239E339",
		x"E439E539", x"E639E739", x"E839E939", x"EA39EB39", x"EC39ED39", x"EE39EF39", x"F039F139", x"F239F339",
		x"F439F539", x"F639F739", x"F839F939", x"FA39FB39", x"FC39FD39", x"FE39FF39", x"FFFFFFFF", x"FFFFFFFF",
		x"003A013A", x"023A033A", x"043A053A", x"063A073A", x"083A093A", x"0A3A0B3A", x"0C3A0D3A", x"0E3A0F3A",
		x"103A113A", x"123A133A", x"143A153A", x"163A173A", x"183A193A", x"1A3A1B3A", x"1C3A1D3A", x"1E3A1F3A",
		x"203A213A", x"223A233A", x"243A253A", x"263A273A", x"283A293A", x"2A3A2B3A", x"2C3A2D3A", x"2E3A2F3A",
		x"303A313A", x"323A333A", x"343A353A", x"363A373A", x"383A393A", x"3A3A3B3A", x"3C3A3D3A", x"3E3A3F3A",
		x"FFFFFFFF", x"FFFFFFFF", x"403A413A", x"423A433A", x"443A453A", x"463A473A", x"483A493A", x"4A3A4B3A",
		x"4C3A4D3A", x"4E3A4F3A", x"503A513A", x"523A533A", x"543A553A", x"563A573A", x"583A593A", x"5A3A5B3A",
		x"5C3A5D3A", x"5E3A5F3A", x"603A613A", x"623A633A", x"643A653A", x"663A673A", x"683A693A", x"6A3A6B3A",
		x"6C3A6D3A", x"6E3A6F3A", x"703A713A", x"723A733A", x"743A753A", x"763A773A", x"783A793A", x"7A3A7B3A",
		x"7C3A7D3A", x"7E3A7F3A", x"FFFFFFFF", x"FFFFFFFF", x"803A813A", x"823A833A", x"843A853A", x"863A873A",
		x"883A893A", x"8A3A8B3A", x"8C3A8D3A", x"8E3A8F3A", x"903A913A", x"923A933A", x"943A953A", x"963A973A",
		x"983A993A", x"9A3A9B3A", x"9C3A9D3A", x"9E3A9F3A", x"A03AA13A", x"A23AA33A", x"A43AA53A", x"A63AA73A",
		x"A83AA93A", x"AA3AAB3A", x"AC3AAD3A", x"AE3AAF3A", x"B03AB13A", x"B23AB33A", x"B43AB53A", x"B63AB73A",
		x"B83AB93A", x"BA3ABB3A", x"BC3ABD3A", x"BE3ABF3A", x"FFFFFFFF", x"FFFFFFFF", x"C03AC13A", x"C23AC33A",
		x"C43AC53A", x"C63AC73A", x"C83AC93A", x"CA3ACB3A", x"CC3ACD3A", x"CE3ACF3A", x"D03AD13A", x"D23AD33A",
		x"D43AD53A", x"D63AD73A", x"D83AD93A", x"DA3ADB3A", x"DC3ADD3A", x"DE3ADF3A", x"E03AE13A", x"E23AE33A",
		x"E43AE53A", x"E63AE73A", x"E83AE93A", x"EA3AEB3A", x"EC3AED3A", x"EE3AEF3A", x"F03AF13A", x"F23AF33A",
		x"F43AF53A", x"F63AF73A", x"F83AF93A", x"FA3AFB3A", x"FC3AFD3A", x"FE3AFF3A", x"FFFFFFFF", x"FFFFFFFF",
		x"003B013B", x"023B033B", x"043B053B", x"063B073B", x"083B093B", x"0A3B0B3B", x"0C3B0D3B", x"0E3B0F3B",
		x"103B113B", x"123B133B", x"143B153B", x"163B173B", x"183B193B", x"1A3B1B3B", x"1C3B1D3B", x"1E3B1F3B",
		x"203B213B", x"223B233B", x"243B253B", x"263B273B", x"283B293B", x"2A3B2B3B", x"2C3B2D3B", x"2E3B2F3B",
		x"303B313B", x"323B333B", x"343B353B", x"363B373B", x"383B393B", x"3A3B3B3B", x"3C3B3D3B", x"3E3B3F3B",
		x"FFFFFFFF", x"FFFFFFFF", x"403B413B", x"423B433B", x"443B453B", x"463B473B", x"483B493B", x"4A3B4B3B",
		x"4C3B4D3B", x"4E3B4F3B", x"503B513B", x"523B533B", x"543B553B", x"563B573B", x"583B593B", x"5A3B5B3B",
		x"5C3B5D3B", x"5E3B5F3B", x"603B613B", x"623B633B", x"643B653B", x"663B673B", x"683B693B", x"6A3B6B3B",
		x"6C3B6D3B", x"6E3B6F3B", x"703B713B", x"723B733B", x"743B753B", x"763B773B", x"783B793B", x"7A3B7B3B",
		x"7C3B7D3B", x"7E3B7F3B", x"FFFFFFFF", x"FFFFFFFF", x"803B813B", x"823B833B", x"843B853B", x"863B873B",
		x"883B893B", x"8A3B8B3B", x"8C3B8D3B", x"8E3B8F3B", x"903B913B", x"923B933B", x"943B953B", x"963B973B",
		x"983B993B", x"9A3B9B3B", x"9C3B9D3B", x"9E3B9F3B", x"A03BA13B", x"A23BA33B", x"A43BA53B", x"A63BA73B",
		x"A83BA93B", x"AA3BAB3B", x"AC3BAD3B", x"AE3BAF3B", x"B03BB13B", x"B23BB33B", x"B43BB53B", x"B63BB73B",
		x"B83BB93B", x"BA3BBB3B", x"BC3BBD3B", x"BE3BBF3B", x"FFFFFFFF", x"FFFFFFFF", x"C03BC13B", x"C23BC33B",
		x"C43BC53B", x"C63BC73B", x"C83BC93B", x"CA3BCB3B", x"CC3BCD3B", x"CE3BCF3B", x"D03BD13B", x"D23BD33B",
		x"D43BD53B", x"D63BD73B", x"D83BD93B", x"DA3BDB3B", x"DC3BDD3B", x"DE3BDF3B", x"E03BE13B", x"E23BE33B",
		x"E43BE53B", x"E63BE73B", x"E83BE93B", x"EA3BEB3B", x"EC3BED3B", x"EE3BEF3B", x"F03BF13B", x"F23BF33B",
		x"F43BF53B", x"F63BF73B", x"F83BF93B", x"FA3BFB3B", x"FC3BFD3B", x"FE3BFF3B", x"FFFFFFFF", x"FFFFFFFF",
		x"003C013C", x"023C033C", x"043C053C", x"063C073C", x"083C093C", x"0A3C0B3C", x"0C3C0D3C", x"0E3C0F3C",
		x"103C113C", x"123C133C", x"143C153C", x"163C173C", x"183C193C", x"1A3C1B3C", x"1C3C1D3C", x"1E3C1F3C",
		x"203C213C", x"223C233C", x"243C253C", x"263C273C", x"283C293C", x"2A3C2B3C", x"2C3C2D3C", x"2E3C2F3C",
		x"303C313C", x"323C333C", x"343C353C", x"363C373C", x"383C393C", x"3A3C3B3C", x"3C3C3D3C", x"3E3C3F3C",
		x"FFFFFFFF", x"FFFFFFFF", x"403C413C", x"423C433C", x"443C453C", x"463C473C", x"483C493C", x"4A3C4B3C",
		x"4C3C4D3C", x"4E3C4F3C", x"503C513C", x"523C533C", x"543C553C", x"563C573C", x"583C593C", x"5A3C5B3C",
		x"5C3C5D3C", x"5E3C5F3C", x"603C613C", x"623C633C", x"643C653C", x"663C673C", x"683C693C", x"6A3C6B3C",
		x"6C3C6D3C", x"6E3C6F3C", x"703C713C", x"723C733C", x"743C753C", x"763C773C", x"783C793C", x"7A3C7B3C",
		x"7C3C7D3C", x"7E3C7F3C", x"FFFFFFFF", x"FFFFFFFF", x"803C813C", x"823C833C", x"843C853C", x"863C873C",
		x"883C893C", x"8A3C8B3C", x"8C3C8D3C", x"8E3C8F3C", x"903C913C", x"923C933C", x"943C953C", x"963C973C",
		x"983C993C", x"9A3C9B3C", x"9C3C9D3C", x"9E3C9F3C", x"A03CA13C", x"A23CA33C", x"A43CA53C", x"A63CA73C",
		x"A83CA93C", x"AA3CAB3C", x"AC3CAD3C", x"AE3CAF3C", x"B03CB13C", x"B23CB33C", x"B43CB53C", x"B63CB73C",
		x"B83CB93C", x"BA3CBB3C", x"BC3CBD3C", x"BE3CBF3C", x"FFFFFFFF", x"FFFFFFFF", x"C03CC13C", x"C23CC33C",
		x"C43CC53C", x"C63CC73C", x"C83CC93C", x"CA3CCB3C", x"CC3CCD3C", x"CE3CCF3C", x"D03CD13C", x"D23CD33C",
		x"D43CD53C", x"D63CD73C", x"D83CD93C", x"DA3CDB3C", x"DC3CDD3C", x"DE3CDF3C", x"E03CE13C", x"E23CE33C",
		x"E43CE53C", x"E63CE73C", x"E83CE93C", x"EA3CEB3C", x"EC3CED3C", x"EE3CEF3C", x"F03CF13C", x"F23CF33C",
		x"F43CF53C", x"F63CF73C", x"F83CF93C", x"FA3CFB3C", x"FC3CFD3C", x"FE3CFF3C", x"FFFFFFFF", x"FFFFFFFF",
		x"003D013D", x"023D033D", x"043D053D", x"063D073D", x"083D093D", x"0A3D0B3D", x"0C3D0D3D", x"0E3D0F3D",
		x"103D113D", x"123D133D", x"143D153D", x"163D173D", x"183D193D", x"1A3D1B3D", x"1C3D1D3D", x"1E3D1F3D",
		x"203D213D", x"223D233D", x"243D253D", x"263D273D", x"283D293D", x"2A3D2B3D", x"2C3D2D3D", x"2E3D2F3D",
		x"303D313D", x"323D333D", x"343D353D", x"363D373D", x"383D393D", x"3A3D3B3D", x"3C3D3D3D", x"3E3D3F3D",
		x"FFFFFFFF", x"FFFFFFFF", x"403D413D", x"423D433D", x"443D453D", x"463D473D", x"483D493D", x"4A3D4B3D",
		x"4C3D4D3D", x"4E3D4F3D", x"503D513D", x"523D533D", x"543D553D", x"563D573D", x"583D593D", x"5A3D5B3D",
		x"5C3D5D3D", x"5E3D5F3D", x"603D613D", x"623D633D", x"643D653D", x"663D673D", x"683D693D", x"6A3D6B3D",
		x"6C3D6D3D", x"6E3D6F3D", x"703D713D", x"723D733D", x"743D753D", x"763D773D", x"783D793D", x"7A3D7B3D",
		x"7C3D7D3D", x"7E3D7F3D", x"FFFFFFFF", x"FFFFFFFF", x"803D813D", x"823D833D", x"843D853D", x"863D873D",
		x"883D893D", x"8A3D8B3D", x"8C3D8D3D", x"8E3D8F3D", x"903D913D", x"923D933D", x"943D953D", x"963D973D",
		x"983D993D", x"9A3D9B3D", x"9C3D9D3D", x"9E3D9F3D", x"A03DA13D", x"A23DA33D", x"A43DA53D", x"A63DA73D",
		x"A83DA93D", x"AA3DAB3D", x"AC3DAD3D", x"AE3DAF3D", x"B03DB13D", x"B23DB33D", x"B43DB53D", x"B63DB73D",
		x"B83DB93D", x"BA3DBB3D", x"BC3DBD3D", x"BE3DBF3D", x"FFFFFFFF", x"FFFFFFFF", x"C03DC13D", x"C23DC33D",
		x"C43DC53D", x"C63DC73D", x"C83DC93D", x"CA3DCB3D", x"CC3DCD3D", x"CE3DCF3D", x"D03DD13D", x"D23DD33D",
		x"D43DD53D", x"D63DD73D", x"D83DD93D", x"DA3DDB3D", x"DC3DDD3D", x"DE3DDF3D", x"E03DE13D", x"E23DE33D",
		x"E43DE53D", x"E63DE73D", x"E83DE93D", x"EA3DEB3D", x"EC3DED3D", x"EE3DEF3D", x"F03DF13D", x"F23DF33D",
		x"F43DF53D", x"F63DF73D", x"F83DF93D", x"FA3DFB3D", x"FC3DFD3D", x"FE3DFF3D", x"FFFFFFFF", x"FFFFFFFF",
		x"003E013E", x"023E033E", x"043E053E", x"063E073E", x"083E093E", x"0A3E0B3E", x"0C3E0D3E", x"0E3E0F3E",
		x"103E113E", x"123E133E", x"143E153E", x"163E173E", x"183E193E", x"1A3E1B3E", x"1C3E1D3E", x"1E3E1F3E",
		x"203E213E", x"223E233E", x"243E253E", x"263E273E", x"283E293E", x"2A3E2B3E", x"2C3E2D3E", x"2E3E2F3E",
		x"303E313E", x"323E333E", x"343E353E", x"363E373E", x"383E393E", x"3A3E3B3E", x"3C3E3D3E", x"3E3E3F3E",
		x"FFFFFFFF", x"FFFFFFFF", x"403E413E", x"423E433E", x"443E453E", x"463E473E", x"483E493E", x"4A3E4B3E",
		x"4C3E4D3E", x"4E3E4F3E", x"503E513E", x"523E533E", x"543E553E", x"563E573E", x"583E593E", x"5A3E5B3E",
		x"5C3E5D3E", x"5E3E5F3E", x"603E613E", x"623E633E", x"643E653E", x"663E673E", x"683E693E", x"6A3E6B3E",
		x"6C3E6D3E", x"6E3E6F3E", x"703E713E", x"723E733E", x"743E753E", x"763E773E", x"783E793E", x"7A3E7B3E",
		x"7C3E7D3E", x"7E3E7F3E", x"FFFFFFFF", x"FFFFFFFF", x"803E813E", x"823E833E", x"843E853E", x"863E873E",
		x"883E893E", x"8A3E8B3E", x"8C3E8D3E", x"8E3E8F3E", x"903E913E", x"923E933E", x"943E953E", x"963E973E",
		x"983E993E", x"9A3E9B3E", x"9C3E9D3E", x"9E3E9F3E", x"A03EA13E", x"A23EA33E", x"A43EA53E", x"A63EA73E",
		x"A83EA93E", x"AA3EAB3E", x"AC3EAD3E", x"AE3EAF3E", x"B03EB13E", x"B23EB33E", x"B43EB53E", x"B63EB73E",
		x"B83EB93E", x"BA3EBB3E", x"BC3EBD3E", x"BE3EBF3E", x"FFFFFFFF", x"FFFFFFFF", x"C03EC13E", x"C23EC33E",
		x"C43EC53E", x"C63EC73E", x"C83EC93E", x"CA3ECB3E", x"CC3ECD3E", x"CE3ECF3E", x"D03ED13E", x"D23ED33E",
		x"D43ED53E", x"D63ED73E", x"D83ED93E", x"DA3EDB3E", x"DC3EDD3E", x"DE3EDF3E", x"E03EE13E", x"E23EE33E",
		x"E43EE53E", x"E63EE73E", x"E83EE93E", x"EA3EEB3E", x"EC3EED3E", x"EE3EEF3E", x"F03EF13E", x"F23EF33E",
		x"F43EF53E", x"F63EF73E", x"F83EF93E", x"FA3EFB3E", x"FC3EFD3E", x"FE3EFF3E", x"FFFFFFFF", x"FFFFFFFF",
		x"003F013F", x"023F033F", x"043F053F", x"063F073F", x"083F093F", x"0A3F0B3F", x"0C3F0D3F", x"0E3F0F3F",
		x"103F113F", x"123F133F", x"143F153F", x"163F173F", x"183F193F", x"1A3F1B3F", x"1C3F1D3F", x"1E3F1F3F",
		x"203F213F", x"223F233F", x"243F253F", x"263F273F", x"283F293F", x"2A3F2B3F", x"2C3F2D3F", x"2E3F2F3F",
		x"303F313F", x"323F333F", x"343F353F", x"363F373F", x"383F393F", x"3A3F3B3F", x"3C3F3D3F", x"3E3F3F3F",
		x"FFFFFFFF", x"FFFFFFFF", x"403F413F", x"423F433F", x"443F453F", x"463F473F", x"483F493F", x"4A3F4B3F",
		x"4C3F4D3F", x"4E3F4F3F", x"503F513F", x"523F533F", x"543F553F", x"563F573F", x"583F593F", x"5A3F5B3F",
		x"5C3F5D3F", x"5E3F5F3F", x"603F613F", x"623F633F", x"643F653F", x"663F673F", x"683F693F", x"6A3F6B3F",
		x"6C3F6D3F", x"6E3F6F3F", x"703F713F", x"723F733F", x"743F753F", x"763F773F", x"783F793F", x"7A3F7B3F",
		x"7C3F7D3F", x"7E3F7F3F", x"FFFFFFFF", x"FFFFFFFF", x"803F813F", x"823F833F", x"843F853F", x"863F873F",
		x"883F893F", x"8A3F8B3F", x"8C3F8D3F", x"8E3F8F3F", x"903F913F", x"923F933F", x"943F953F", x"963F973F",
		x"983F993F", x"9A3F9B3F", x"9C3F9D3F", x"9E3F9F3F", x"A03FA13F", x"A23FA33F", x"A43FA53F", x"A63FA73F",
		x"A83FA93F", x"AA3FAB3F", x"AC3FAD3F", x"AE3FAF3F", x"B03FB13F", x"B23FB33F", x"B43FB53F", x"B63FB73F",
		x"B83FB93F", x"BA3FBB3F", x"BC3FBD3F", x"BE3FBF3F", x"FFFFFFFF", x"FFFFFFFF", x"C03FC13F", x"C23FC33F",
		x"C43FC53F", x"C63FC73F", x"C83FC93F", x"CA3FCB3F", x"CC3FCD3F", x"CE3FCF3F", x"D03FD13F", x"D23FD33F",
		x"D43FD53F", x"D63FD73F", x"D83FD93F", x"DA3FDB3F", x"DC3FDD3F", x"DE3FDF3F", x"E03FE13F", x"E23FE33F",
		x"E43FE53F", x"E63FE73F", x"E83FE93F", x"EA3FEB3F", x"EC3FED3F", x"EE3FEF3F", x"F03FF13F", x"F23FF33F",
		x"F43FF53F", x"F63FF73F", x"F83FF93F", x"FA3FFB3F", x"FC3FFD3F", x"FE3FFF3F", x"FFFFFFFF", x"FFFFFFFF",
		x"F9602EB1", c_FTDI_PROT_END_OF_PAYLOAD
	);

	-- Imagette Package
	type t_ftdi_prot_imagette_package is array (0 to 7) of std_logic_vector(31 downto 0);
	constant c_FTDI_PROT_IMAGETTE_PACKAGE : t_ftdi_prot_imagette_package := (
		c_FTDI_PROT_START_OF_PACKAGE,
		c_FTDI_PROT_PKG_ID_IMAGETTE_TRANSMISSION,
		x"01020300",
		x"07001000",
		x"6B030000",
		x"00020000",
		x"DC05A26D",
		c_FTDI_PROT_END_OF_HEADER
	);

	-- Imagette Payload
	type t_ftdi_prot_imagette_payload is array (0 to (128 - 1 + 3)) of std_logic_vector(31 downto 0);
	constant c_FTDI_PROT_IMAGETTE_PAYLOAD : t_ftdi_prot_imagette_payload := (
		c_FTDI_PROT_START_OF_PAYLOAD,
		x"11110000", x"33332222", x"55554444", x"77776666", x"99998888", x"BBBBAAAA", x"DDDDCCCC", x"FFFFEEEE",
		x"00000100", x"02000300", x"04000500", x"06000700", x"08000900", x"0A000B00", x"0C000D00", x"0E000F00",
		x"10001100", x"12001300", x"14001500", x"16001700", x"18001900", x"1A001B00", x"1C001D00", x"1E001F00",
		x"20002100", x"22002300", x"24002500", x"26002700", x"28002900", x"2A002B00", x"2C002D00", x"2E002F00",
		x"30003100", x"32003300", x"34003500", x"36003700", x"38003900", x"3A003B00", x"3C003D00", x"3E003F00",
		x"FFFFFFFF", x"FFFFFFFF", x"40004100", x"42004300", x"44004500", x"46004700", x"48004900", x"4A004B00",
		x"4C004D00", x"4E004F00", x"50005100", x"52005300", x"54005500", x"56005700", x"58005900", x"5A005B00",
		x"5C005D00", x"5E005F00", x"60006100", x"62006300", x"64006500", x"66006700", x"68006900", x"6A006B00",
		x"6C006D00", x"6E006F00", x"70007100", x"72007300", x"74007500", x"76007700", x"78007900", x"7A007B00",
		x"7C007D00", x"7E007F00", x"FFFFFFFF", x"FFFFFFFF", x"80008100", x"82008300", x"84008500", x"86008700",
		x"88008900", x"8A008B00", x"8C008D00", x"8E008F00", x"90009100", x"92009300", x"94009500", x"96009700",
		x"98009900", x"9A009B00", x"9C009D00", x"9E009F00", x"A000A100", x"A200A300", x"A400A500", x"A600A700",
		x"A800A900", x"AA00AB00", x"AC00AD00", x"AE00AF00", x"B000B100", x"B200B300", x"B400B500", x"B600B700",
		x"B800B900", x"BA00BB00", x"BC00BD00", x"BE00BF00", x"FFFFFFFF", x"FFFFFFFF", x"C000C100", x"C200C300",
		x"C400C500", x"C600C700", x"C800C900", x"CA00CB00", x"CC00CD00", x"CE00CF00", x"D000D100", x"D200D300",
		x"D400D500", x"D600D700", x"D800D900", x"DA00DB00", x"DC00DD00", x"DE00DF00", x"E000E100", x"E200E300",
		x"0F9C40BB", c_FTDI_PROT_END_OF_PAYLOAD
	);

begin

	-- bidir io buffer instantiation, for the umft601a module pins (fpga <--> umft601a)
	ftdi_inout_io_buffer_39b_inst : entity work.ftdi_inout_io_buffer_39b
		port map(
			datain(38 downto 7)  => s_umft601a_data_out,
			datain(6)            => s_umft601a_wakeup_n_out,
			datain(5 downto 2)   => s_umft601a_be_out,
			datain(1 downto 0)   => s_umft601a_gpio_out,
			oe(38)               => s_umft601a_oe,
			oe(37)               => s_umft601a_oe,
			oe(36)               => s_umft601a_oe,
			oe(35)               => s_umft601a_oe,
			oe(34)               => s_umft601a_oe,
			oe(33)               => s_umft601a_oe,
			oe(32)               => s_umft601a_oe,
			oe(31)               => s_umft601a_oe,
			oe(30)               => s_umft601a_oe,
			oe(29)               => s_umft601a_oe,
			oe(28)               => s_umft601a_oe,
			oe(27)               => s_umft601a_oe,
			oe(26)               => s_umft601a_oe,
			oe(25)               => s_umft601a_oe,
			oe(24)               => s_umft601a_oe,
			oe(23)               => s_umft601a_oe,
			oe(22)               => s_umft601a_oe,
			oe(21)               => s_umft601a_oe,
			oe(20)               => s_umft601a_oe,
			oe(19)               => s_umft601a_oe,
			oe(18)               => s_umft601a_oe,
			oe(17)               => s_umft601a_oe,
			oe(16)               => s_umft601a_oe,
			oe(15)               => s_umft601a_oe,
			oe(14)               => s_umft601a_oe,
			oe(13)               => s_umft601a_oe,
			oe(12)               => s_umft601a_oe,
			oe(11)               => s_umft601a_oe,
			oe(10)               => s_umft601a_oe,
			oe(9)                => s_umft601a_oe,
			oe(8)                => s_umft601a_oe,
			oe(7)                => s_umft601a_oe,
			oe(6)                => s_umft601a_oe,
			oe(5)                => s_umft601a_oe,
			oe(4)                => s_umft601a_oe,
			oe(3)                => s_umft601a_oe,
			oe(2)                => s_umft601a_oe,
			oe(1)                => s_umft601a_oe,
			oe(0)                => s_umft601a_oe,
			dataio(38 downto 7)  => umft_data_bus_io,
			dataio(6)            => umft_wakeup_n_pin_io,
			dataio(5 downto 2)   => umft_be_bus_io,
			dataio(1 downto 0)   => umft_gpio_bus_io,
			dataout(38 downto 7) => s_umft601a_data_in,
			dataout(6)           => s_umft601a_wakeup_n_in,
			dataout(5 downto 2)  => s_umft601a_be_in,
			dataout(1 downto 0)  => s_umft601a_gpio_in
		);
	s_umft601a_oe <= not (umft_oe_n_pin_i);

	p_usb3_fifo_master_stimuli : process(clk_i, rst_i) is
		variable v_data_cnt : natural := 0;
	begin
		if (rst_i = '1') then

			umft_rxf_n_pin_o        <= '1';
			umft_txe_n_pin_o        <= '1';
			s_umft601a_data_out     <= (others => '0');
			s_umft601a_wakeup_n_out <= '1';
			s_umft601a_be_out       <= (others => '0');
			s_umft601a_gpio_out     <= (others => '1');
			s_counter               <= 0;
			s_counter2              <= 0;
			v_data_cnt              := 0;
			s_times_cnt             <= 0;

		elsif rising_edge(clk_i) then

			umft_rxf_n_pin_o        <= '1';
			umft_txe_n_pin_o        <= '1';
			s_umft601a_data_out     <= (others => '0');
			s_umft601a_wakeup_n_out <= '1';
			s_umft601a_be_out       <= (others => '0');
			s_umft601a_gpio_out     <= (others => '1');
			s_counter               <= s_counter + 1;
			--			s_counter2              <= s_counter2 + 1;

			case s_counter is
				
-- Imagette Transmission --

				when (33 - 4) to (33 - 1) =>
					umft_rxf_n_pin_o        <= '0';
					umft_txe_n_pin_o        <= '1';
					s_umft601a_data_out     <= (others => '0');
					s_umft601a_wakeup_n_out <= '1';
					s_umft601a_be_out       <= (others => '0');
					s_umft601a_gpio_out     <= (others => '1');
					v_data_cnt              := 0;

				when 33 to (33 - 1 + 8) =>
					umft_rxf_n_pin_o        <= '0';
					umft_txe_n_pin_o        <= '1';
					s_umft601a_data_out     <= c_FTDI_PROT_IMAGETTE_PACKAGE(v_data_cnt);
					v_data_cnt              := v_data_cnt + 1;
					s_umft601a_wakeup_n_out <= '1';
					s_umft601a_be_out       <= (others => '1');
					s_umft601a_gpio_out     <= (others => '1');

				when (33 + 8) =>
					umft_rxf_n_pin_o        <= '1';
					umft_txe_n_pin_o        <= '1';
					s_umft601a_data_out     <= (others => '0');
					s_umft601a_wakeup_n_out <= '1';
					s_umft601a_be_out       <= (others => '0');
					s_umft601a_gpio_out     <= (others => '1');
					v_data_cnt              := 0;

				when (100 - 4) to (100 - 1) =>
					umft_rxf_n_pin_o        <= '0';
					umft_txe_n_pin_o        <= '1';
					s_umft601a_data_out     <= (others => '0');
					s_umft601a_wakeup_n_out <= '1';
					s_umft601a_be_out       <= (others => '0');
					s_umft601a_gpio_out     <= (others => '1');
					v_data_cnt              := 0;

								when 100 to (100 - 1 + 1024) =>
				--					if (umft_rd_n_pin_i = '0') then
										umft_rxf_n_pin_o        <= '0';
										umft_txe_n_pin_o        <= '1';
										if (v_data_cnt < (t_ftdi_prot_imagette_payload'high + 1)) then
											s_umft601a_data_out     <= c_FTDI_PROT_IMAGETTE_PAYLOAD(v_data_cnt);
										else
											s_umft601a_data_out     <= (others => '0');
										end if;
										v_data_cnt              := v_data_cnt + 1;
										s_umft601a_wakeup_n_out <= '1';
										s_umft601a_be_out       <= (others => '1');
										s_umft601a_gpio_out     <= (others => '1');
				--					else
				--						umft_rxf_n_pin_o        <= '0';
				--						umft_txe_n_pin_o        <= '1';
				--						s_umft601a_data_out     <= (others => '0');
				--						s_umft601a_wakeup_n_out <= '1';
				--						s_umft601a_be_out       <= (others => '1');
				--						s_umft601a_gpio_out     <= (others => '1');
				--						s_counter               <= s_counter;
				--					end if;
					
								when (100 + 1024) =>
									umft_rxf_n_pin_o        <= '1';
									umft_txe_n_pin_o        <= '1';
									s_umft601a_data_out     <= (others => '0');
									s_umft601a_wakeup_n_out <= '1';
									s_umft601a_be_out       <= (others => '0');
									s_umft601a_gpio_out     <= (others => '1');
										if (s_counter = (100 + 1024)) then
											if (s_counter2 = 10) then
												s_counter  <= 10000;
												s_counter2 <= 0;
												v_data_cnt              := 0;
											else
												s_counter  <= 1000;
												s_counter2 <= s_counter2 + 1;
											end if;
										end if;

				---------------------------
				
				---- LUT Transmission -----

--				when (33 - 4) to (33 - 1) =>
--					umft_rxf_n_pin_o        <= '0';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= (others => '0');
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '0');
--					s_umft601a_gpio_out     <= (others => '1');
--					v_data_cnt              := 0;
--
--				when 33 to (33 - 1 + 8) =>
--					umft_rxf_n_pin_o        <= '0';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= c_FTDI_PROT_ACK_PACKAGE(v_data_cnt);
--					v_data_cnt              := v_data_cnt + 1;
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '1');
--					s_umft601a_gpio_out     <= (others => '1');
--
--				when (33 + 8) =>
--					umft_rxf_n_pin_o        <= '1';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= (others => '0');
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '0');
--					s_umft601a_gpio_out     <= (others => '1');
--					v_data_cnt              := 0;
--
--				when (400 - 4) to (400 - 1) =>
--					umft_rxf_n_pin_o        <= '0';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= (others => '0');
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '0');
--					s_umft601a_gpio_out     <= (others => '1');
--					v_data_cnt              := 0;
--
--				when 400 to (400 - 1 + 8) =>
--					umft_rxf_n_pin_o        <= '0';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= c_FTDI_PROT_ACK_PACKAGE(v_data_cnt);
--					v_data_cnt              := v_data_cnt + 1;
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '1');
--					s_umft601a_gpio_out     <= (others => '1');
--
--				when (400 + 8) =>
--					umft_rxf_n_pin_o        <= '1';
--					umft_txe_n_pin_o        <= '1';
--					s_umft601a_data_out     <= (others => '0');
--					s_umft601a_wakeup_n_out <= '1';
--					s_umft601a_be_out       <= (others => '0');
--					s_umft601a_gpio_out     <= (others => '1');
--					v_data_cnt              := 0;
					
					---------------------------
					
					--- Full-Image Request ----

				--				when 69 to 72 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--
				--				when 73 to (73 - 1 + 8) =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= c_FTDI_PROT_REPLY_PACKAGE(v_data_cnt);
				--					v_data_cnt              := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '1');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					
				--				when (73 + 8) =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--					s_counter               <= 5000;
				--
				--				when 5099 to 5102 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--
				--				when 5103 to (5103 - 1 + 1024) =>
				----					if (umft_rd_n_pin_i = '0') then
				--						umft_rxf_n_pin_o        <= '0';
				--						umft_txe_n_pin_o        <= '1';
				--						if (v_data_cnt < (t_ftdi_prot_reply_payload'high + 1)) then
				--							s_umft601a_data_out     <= c_FTDI_PROT_REPLY_PAYLOAD(v_data_cnt);
				--						else
				--							s_umft601a_data_out     <= (others => '0');
				--						end if;
				--						v_data_cnt              := v_data_cnt + 1;
				--						s_umft601a_wakeup_n_out <= '1';
				--						s_umft601a_be_out       <= (others => '1');
				--						s_umft601a_gpio_out     <= (others => '1');
				----					else
				----						umft_rxf_n_pin_o        <= '0';
				----						umft_txe_n_pin_o        <= '1';
				----						s_umft601a_data_out     <= (others => '0');
				----						s_umft601a_wakeup_n_out <= '1';
				----						s_umft601a_be_out       <= (others => '1');
				----						s_umft601a_gpio_out     <= (others => '1');
				----						s_counter               <= s_counter;
				----					end if;
				--
				--				when (5103 + 1024) =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--						if (s_counter = (5103 + 1024)) then
				--							if (s_counter2 = 10) then
				--								s_counter  <= 10000;
				--								s_counter2 <= 0;
				--								v_data_cnt              := 0;
				--							else
				--								s_counter  <= 1000;
				--								s_counter2 <= s_counter2 + 1;
				--							end if;
				--						end if;

				--												when 10000 to 10002 =>
				--													umft_rxf_n_pin_o        <= '0';
				--													umft_txe_n_pin_o        <= '1';
				--													s_umft601a_data_out     <= (others => '0');
				--													s_umft601a_wakeup_n_out <= '1';
				--													s_umft601a_be_out       <= (others => '0');
				--													s_umft601a_gpio_out     <= (others => '1');
				--													v_data_cnt              := 0;
				--								
				--												when 10003 to (10003 - 1 + 1024) =>
				--													umft_rxf_n_pin_o                  <= '0';
				--													umft_txe_n_pin_o                  <= '1';
				--													s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--													v_data_cnt                        := v_data_cnt + 1;
				--													s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--													v_data_cnt                        := v_data_cnt + 1;
				--													s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--													v_data_cnt                        := v_data_cnt + 1;
				--													s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--													v_data_cnt                        := v_data_cnt + 1;
				--													s_umft601a_wakeup_n_out           <= '1';
				--													s_umft601a_be_out                 <= (others => '1');
				--													s_umft601a_gpio_out               <= (others => '1');
				
				---------------------------
				
				--
				--				when (2503 + 1024) =>
				--					if (s_times_cnt >= (8 - 1)) then
				--						s_times_cnt <= 0;
				--					else
				--						s_times_cnt <= s_times_cnt + 1;
				--						s_counter   <= 2500 - 2000;
				--					end if;

				--				when 3500 to 3502 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--				
				--				when 3503 to (3503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o                  <= '0';
				--					umft_txe_n_pin_o                  <= '1';
				--					s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out           <= '1';
				--					s_umft601a_be_out                 <= (others => '1');
				--					s_umft601a_gpio_out               <= (others => '1');
				--					
				--				when 5500 to 5502 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--					
				--				when 5503 to (5503 - 1 + 512) =>
				--					umft_rxf_n_pin_o                  <= '0';
				--					umft_txe_n_pin_o                  <= '1';
				--					s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out           <= '1';
				--					s_umft601a_be_out                 <= (others => '1');
				--					s_umft601a_gpio_out               <= (others => '1');
				--					
				--				when 7500 to 7502 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--					
				--				when 7503 to (7503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o                  <= '0';
				--					umft_txe_n_pin_o                  <= '1';
				--					s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out           <= '1';
				--					s_umft601a_be_out                 <= (others => '1');
				--					s_umft601a_gpio_out               <= (others => '1');
				--					
				--				when 9500 to 9502 =>
				--					umft_rxf_n_pin_o        <= '0';
				--					umft_txe_n_pin_o        <= '1';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--					
				--				when 9503 to (9503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o                  <= '0';
				--					umft_txe_n_pin_o                  <= '1';
				--					s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out           <= '1';
				--					s_umft601a_be_out                 <= (others => '1');
				--					s_umft601a_gpio_out               <= (others => '1');

				--				when (1503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o                  <= '0';
				--					umft_txe_n_pin_o                  <= '1';
				--					s_umft601a_data_out(31 downto 24) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(23 downto 16) <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(15 downto 8)  <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_data_out(7 downto 0)   <= std_logic_vector(to_unsigned(v_data_cnt, 8));
				--					v_data_cnt                        := v_data_cnt + 1;
				--					s_umft601a_wakeup_n_out           <= '1';
				--					s_umft601a_be_out(3)               <= '0';
				--					s_umft601a_be_out(2)               <= '0';
				--					s_umft601a_be_out(1)               <= '0';
				--					s_umft601a_be_out(0)               <= '1';
				--					s_umft601a_gpio_out               <= (others => '1');

				--												when 60000 to 60002 =>
				--													umft_rxf_n_pin_o        <= '1';
				--													umft_txe_n_pin_o        <= '0';
				--													s_umft601a_data_out     <= (others => '0');
				--													s_umft601a_wakeup_n_out <= '1';
				--													s_umft601a_be_out       <= (others => '0');
				--													s_umft601a_gpio_out     <= (others => '1');
				--													v_data_cnt              := 0;
				--								
				--												when 60003 to (60003 - 1 + 1024) =>
				--													umft_rxf_n_pin_o        <= '1';
				--													umft_txe_n_pin_o        <= '0';
				--													s_umft601a_data_out     <= (others => '0');
				--													s_umft601a_wakeup_n_out <= '1';
				--													s_umft601a_be_out       <= (others => '0');
				--													s_umft601a_gpio_out     <= (others => '1');
				--													v_data_cnt              := 0;
				--													
				--												when 70000 to 70002 =>
				--													umft_rxf_n_pin_o        <= '1';
				--													umft_txe_n_pin_o        <= '0';
				--													s_umft601a_data_out     <= (others => '0');
				--													s_umft601a_wakeup_n_out <= '1';
				--													s_umft601a_be_out       <= (others => '0');
				--													s_umft601a_gpio_out     <= (others => '1');
				--													v_data_cnt              := 0;
				--								
				--												when 70003 to (70003 - 1 + 1024) =>
				--													umft_rxf_n_pin_o        <= '1';
				--													umft_txe_n_pin_o        <= '0';
				--													s_umft601a_data_out     <= (others => '0');
				--													s_umft601a_wakeup_n_out <= '1';
				--													s_umft601a_be_out       <= (others => '0');
				--													s_umft601a_gpio_out     <= (others => '1');
				--													v_data_cnt              := 0;

				--				when (60003 + 1024) =>
				--					if (s_times_cnt >= (8 - 1)) then
				--						s_times_cnt <= 0;
				--					else
				--						s_times_cnt <= s_times_cnt + 1;
				--						s_counter   <= 60000 - 2000;
				--					end if;
				--					
				--				when 2500 to 2502 =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '0';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--
				--				when 2503 to (2503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '0';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;

				--								when 3500 to 3502 =>
				--									umft_rxf_n_pin_o        <= '1';
				--									umft_txe_n_pin_o        <= '0';
				--									s_umft601a_data_out     <= (others => '0');
				--									s_umft601a_wakeup_n_out <= '1';
				--									s_umft601a_be_out       <= (others => '0');
				--									s_umft601a_gpio_out     <= (others => '1');
				--									v_data_cnt              := 0;
				--				
				--								when 3503 to (3503 - 1 + 6) =>
				--									umft_rxf_n_pin_o        <= '1';
				--									umft_txe_n_pin_o        <= '0';
				--									s_umft601a_data_out     <= (others => '0');
				--									s_umft601a_wakeup_n_out <= '1';
				--									s_umft601a_be_out       <= (others => '0');
				--									s_umft601a_gpio_out     <= (others => '1');
				--									v_data_cnt              := 0;
				--					
				--				when 15500 to 15502 =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '0';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;
				--
				--				when 15503 to (15503 - 1 + 1024) =>
				--					umft_rxf_n_pin_o        <= '1';
				--					umft_txe_n_pin_o        <= '0';
				--					s_umft601a_data_out     <= (others => '0');
				--					s_umft601a_wakeup_n_out <= '1';
				--					s_umft601a_be_out       <= (others => '0');
				--					s_umft601a_gpio_out     <= (others => '1');
				--					v_data_cnt              := 0;

				--				when 15000 =>
				--					s_counter               <= 0;

				when others =>
					null;

			end case;

			--			umft_txe_n_pin_o        <= '1';
			--			
			--			case s_counter2 is
			--				
			--				when 2526 to 2528 =>
			--					umft_txe_n_pin_o        <= '0';
			--
			--				when 2529 to (2529 - 1 + 1024) =>
			--					umft_txe_n_pin_o        <= '0';
			--					
			--				when others =>
			--					null;
			--
			--			end case;

		end if;
	end process p_usb3_fifo_master_stimuli;

end architecture RTL;
