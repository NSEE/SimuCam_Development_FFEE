RX_LVDS_inst : RX_LVDS PORT MAP (
		rx_in	 => rx_in_sig,
		rx_out	 => rx_out_sig
	);
