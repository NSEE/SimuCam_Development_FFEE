ftdi_inout_io_buffer_39b_inst : ftdi_inout_io_buffer_39b PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataio	 => dataio_sig,
		dataout	 => dataout_sig
	);
