ftdi_in_io_buffer_3b_inst : ftdi_in_io_buffer_3b PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
