library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity comm_tb_avs_left_read_stimuli is
	generic(
		g_ADDRESS_WIDTH : natural range 1 to 64;
		g_DATA_WIDTH    : natural range 1 to 256
	);
	port(
		clk_i                       : in  std_logic;
		rst_i                       : in  std_logic;
		avs_avalon_mm_address_i     : in  std_logic_vector((g_ADDRESS_WIDTH - 1) downto 0); -- avs_avalon_mm.address
		avs_avalon_mm_read_i        : in  std_logic; --                                     --              .read
		avs_avalon_mm_readata_o     : out std_logic_vector((g_DATA_WIDTH - 1) downto 0); -- --              .readdata
		avs_avalon_mm_waitrequest_o : out std_logic ---                                     --              .waitrequest
	);
end entity comm_tb_avs_left_read_stimuli;

architecture RTL of comm_tb_avs_left_read_stimuli is

	constant c_CCD_IMGDATA_SELECTION : std_logic := '1'; -- '0' = No Data / '1' = With Data

	-- ccd image data
	constant c_CCD_IMGDATA_LENGTH    : natural                                       := 85;
	signal s_ccd_imgdata_cnt         : natural range 0 to (c_CCD_IMGDATA_LENGTH - 1) := 0;
	type t_ccd_imgdata is array (0 to (c_CCD_IMGDATA_LENGTH - 1)) of std_logic_vector(255 downto 0);
	constant c_CCD_IMGDATA_NO_DATA   : t_ccd_imgdata                                 := (
		x"0010000F000E000D000C000B000A000900080007000600050004000300020001",
		x"0020001F001E001D001C001B001A001900180017001600150014001300120011",
		x"0030002F002E002D002C002B002A002900280027002600250024002300220021",
		x"0040003F003E003D003C003B003A003900380037003600350034003300320031",
		x"004C004B004A0049004800470046004500440043004200410000000000000000",
		x"005C005B005A0059005800570056005500540053005200510050004F004E004D",
		x"006C006B006A0069006800670066006500640063006200610060005F005E005D",
		x"007C007B007A0079007800770076007500740073007200710070006F006E006D",
		x"0088008700860085008400830082008100000000000000000080007F007E007D",
		x"009800970096009500940093009200910090008F008E008D008C008B008A0089",
		x"00A800A700A600A500A400A300A200A100A0009F009E009D009C009B009A0099",
		x"00B800B700B600B500B400B300B200B100B000AF00AE00AD00AC00AB00AA00A9",
		x"00C400C300C200C1000000000000000000C000BF00BE00BD00BC00BB00BA00B9",
		x"00D400D300D200D100D000CF00CE00CD00CC00CB00CA00C900C800C700C600C5",
		x"00E400E300E200E100E000DF00DE00DD00DC00DB00DA00D900D800D700D600D5",
		x"00F400F300F200F100F000EF00EE00ED00EC00EB00EA00E900E800E700E600E5",
		x"0000000000000000010000FF00FE00FD00FC00FB00FA00F900F800F700F600F5",
		x"0110010F010E010D010C010B010A010901080107010601050104010301020101",
		x"0120011F011E011D011C011B011A011901180117011601150114011301120111",
		x"0130012F012E012D012C012B012A012901280127012601250124012301220121",
		x"0140013F013E013D013C013B013A013901380137013601350134013301320131",
		x"014C014B014A0149014801470146014501440143014201410000000000000000",
		x"015C015B015A0159015801570156015501540153015201510150014F014E014D",
		x"016C016B016A0169016801670166016501640163016201610160015F015E015D",
		x"017C017B017A0179017801770176017501740173017201710170016F016E016D",
		x"0188018701860185018401830182018100000000000000000180017F017E017D",
		x"019801970196019501940193019201910190018F018E018D018C018B018A0189",
		x"01A801A701A601A501A401A301A201A101A0019F019E019D019C019B019A0199",
		x"01B801B701B601B501B401B301B201B101B001AF01AE01AD01AC01AB01AA01A9",
		x"01C401C301C201C1000000000000000001C001BF01BE01BD01BC01BB01BA01B9",
		x"01D401D301D201D101D001CF01CE01CD01CC01CB01CA01C901C801C701C601C5",
		x"01E401E301E201E101E001DF01DE01DD01DC01DB01DA01D901D801D701D601D5",
		x"01F401F301F201F101F001EF01EE01ED01EC01EB01EA01E901E801E701E601E5",
		x"0000000000000000020001FF01FE01FD01FC01FB01FA01F901F801F701F601F5",
		x"0210020F020E020D020C020B020A020902080207020602050204020302020201",
		x"0220021F021E021D021C021B021A021902180217021602150214021302120211",
		x"0230022F022E022D022C022B022A022902280227022602250224022302220221",
		x"0240023F023E023D023C023B023A023902380237023602350234023302320231",
		x"024C024B024A0249024802470246024502440243024202410000000000000000",
		x"025C025B025A0259025802570256025502540253025202510250024F024E024D",
		x"026C026B026A0269026802670266026502640263026202610260025F025E025D",
		x"027C027B027A0279027802770276027502740273027202710270026F026E026D",
		x"0288028702860285028402830282028100000000000000000280027F027E027D",
		x"029802970296029502940293029202910290028F028E028D028C028B028A0289",
		x"02A802A702A602A502A402A302A202A102A0029F029E029D029C029B029A0299",
		x"02B802B702B602B502B402B302B202B102B002AF02AE02AD02AC02AB02AA02A9",
		x"02C402C302C202C1000000000000000002C002BF02BE02BD02BC02BB02BA02B9",
		x"02D402D302D202D102D002CF02CE02CD02CC02CB02CA02C902C802C702C602C5",
		x"02E402E302E202E102E002DF02DE02DD02DC02DB02DA02D902D802D702D602D5",
		x"02F402F302F202F102F002EF02EE02ED02EC02EB02EA02E902E802E702E602E5",
		x"0000000000000000030002FF02FE02FD02FC02FB02FA02F902F802F702F602F5",
		x"0310030F030E030D030C030B030A030903080307030603050304030303020301",
		x"0320031F031E031D031C031B031A031903180317031603150314031303120311",
		x"0330032F032E032D032C032B032A032903280327032603250324032303220321",
		x"0340033F033E033D033C033B033A033903380337033603350334033303320331",
		x"034C034B034A0349034803470346034503440343034203410000000000000000",
		x"035C035B035A0359035803570356035503540353035203510350034F034E034D",
		x"036C036B036A0369036803670366036503640363036203610360035F035E035D",
		x"037C037B037A0379037803770376037503740373037203710370036F036E036D",
		x"0388038703860385038403830382038100000000000000000380037F037E037D",
		x"039803970396039503940393039203910390038F038E038D038C038B038A0389",
		x"03A803A703A603A503A403A303A203A103A0039F039E039D039C039B039A0399",
		x"03B803B703B603B503B403B303B203B103B003AF03AE03AD03AC03AB03AA03A9",
		x"03C403C303C203C1000000000000000003C003BF03BE03BD03BC03BB03BA03B9",
		x"03D403D303D203D103D003CF03CE03CD03CC03CB03CA03C903C803C703C603C5",
		x"03E403E303E203E103E003DF03DE03DD03DC03DB03DA03D903D803D703D603D5",
		x"03F403F303F203F103F003EF03EE03ED03EC03EB03EA03E903E803E703E603E5",
		x"0000000000000000040003FF03FE03FD03FC03FB03FA03F903F803F703F603F5",
		x"0410040F040E040D040C040B040A040904080407040604050404040304020401",
		x"0420041F041E041D041C041B041A041904180417041604150414041304120411",
		x"0430042F042E042D042C042B042A042904280427042604250424042304220421",
		x"0440043F043E043D043C043B043A043904380437043604350434043304320431",
		x"044C044B044A0449044804470446044504440443044204410000000000000000",
		x"045C045B045A0459045804570456045504540453045204510450044F044E044D",
		x"046C046B046A0469046804670466046504640463046204610460045F045E045D",
		x"047C047B047A0479047804770476047504740473047204710470046F046E046D",
		x"0488048704860485048404830482048100000000000000000480047F047E047D",
		x"049804970496049504940493049204910490048F048E048D048C048B048A0489",
		x"04A804A704A604A504A404A304A204A104A0049F049E049D049C049B049A0499",
		x"04B804B704B604B504B404B304B204B104B004AF04AE04AD04AC04AB04AA04A9",
		x"04C404C304C204C1000000000000000004C004BF04BE04BD04BC04BB04BA04B9",
		x"04D404D304D204D104D004CF04CE04CD04CC04CB04CA04C904C804C704C604C5",
		x"0000000004E204E104E004DF04DE04DD04DC04DB04DA04D904D804D704D604D5",
		x"0000000000000000000000000000000000000000000000000000000000000000",
		x"0000000000000000000000000000000000000000000000000000000000000000"
	);                                  -- no data
	constant c_CCD_IMGDATA_WITH_DATA : t_ccd_imgdata                                 := (
x"0010000F000E000D000C000B000A000900080007000600050004000300020001",
x"0020001F001E001D001C001B001A001900180017001600150014001300120011",
x"0030002F002E002D002C002B002A002900280027002600250024002300220021",
x"0040003F003E003D003C003B003A003900380037003600350034003300320031",
x"004C004B004A004900480047004600450044004300420041FFFFFFFFFFFFFFFF",
x"005C005B005A0059005800570056005500540053005200510050004F004E004D",
x"006C006B006A0069006800670066006500640063006200610060005F005E005D",
x"007C007B007A0079007800770076007500740073007200710070006F006E006D",
x"00880087008600850084008300820081FFFFFFFFFFFFFFFF0080007F007E007D",
x"009800970096009500940093009200910090008F008E008D008C008B008A0089",
x"00A800A700A600A500A400A300A200A100A0009F009E009D009C009B009A0099",
x"00B800B700B600B500B400B300B200B100B000AF00AE00AD00AC00AB00AA00A9",
x"00C400C300C200C1FFFFFFFFFFFFFFFF00C000BF00BE00BD00BC00BB00BA00B9",
x"00D400D300D200D100D000CF00CE00CD00CC00CB00CA00C900C800C700C600C5",
x"00E400E300E200E100E000DF00DE00DD00DC00DB00DA00D900D800D700D600D5",
x"00F400F300F200F100F000EF00EE00ED00EC00EB00EA00E900E800E700E600E5",
x"FFFFFFFFFFFFFFFF010000FF00FE00FD00FC00FB00FA00F900F800F700F600F5",
x"0110010F010E010D010C010B010A010901080107010601050104010301020101",
x"0120011F011E011D011C011B011A011901180117011601150114011301120111",
x"0130012F012E012D012C012B012A012901280127012601250124012301220121",
x"0140013F013E013D013C013B013A013901380137013601350134013301320131",
x"014C014B014A0149014801470146014501440143014201410000000000000000",
x"015C015B015A0159015801570156015501540153015201510150014F014E014D",
x"016C016B016A0169016801670166016501640163016201610160015F015E015D",
x"017C017B017A0179017801770176017501740173017201710170016F016E016D",
x"0188018701860185018401830182018100000000000000000180017F017E017D",
x"019801970196019501940193019201910190018F018E018D018C018B018A0189",
x"01A801A701A601A501A401A301A201A101A0019F019E019D019C019B019A0199",
x"01B801B701B601B501B401B301B201B101B001AF01AE01AD01AC01AB01AA01A9",
x"01C401C301C201C1000000000000000001C001BF01BE01BD01BC01BB01BA01B9",
x"01D401D301D201D101D001CF01CE01CD01CC01CB01CA01C901C801C701C601C5",
x"01E401E301E201E101E001DF01DE01DD01DC01DB01DA01D901D801D701D601D5",
x"01F401F301F201F101F001EF01EE01ED01EC01EB01EA01E901E801E701E601E5",
x"0000000000000000020001FF01FE01FD01FC01FB01FA01F901F801F701F601F5",
x"0210020F020E020D020C020B020A020902080207020602050204020302020201",
x"0220021F021E021D021C021B021A021902180217021602150214021302120211",
x"0230022F022E022D022C022B022A022902280227022602250224022302220221",
x"0240023F023E023D023C023B023A023902380237023602350234023302320231",
x"024C024B024A0249024802470246024502440243024202410000000000000000",
x"025C025B025A0259025802570256025502540253025202510250024F024E024D",
x"026C026B026A0269026802670266026502640263026202610260025F025E025D",
x"027C027B027A0279027802770276027502740273027202710270026F026E026D",
x"0288028702860285028402830282028100000000000000000280027F027E027D",
x"029802970296029502940293029202910290028F028E028D028C028B028A0289",
x"02A802A702A602A502A402A302A202A102A0029F029E029D029C029B029A0299",
x"02B802B702B602B502B402B302B202B102B002AF02AE02AD02AC02AB02AA02A9",
x"02C402C302C202C1000000000000000002C002BF02BE02BD02BC02BB02BA02B9",
x"02D402D302D202D102D002CF02CE02CD02CC02CB02CA02C902C802C702C602C5",
x"02E402E302E202E102E002DF02DE02DD02DC02DB02DA02D902D802D702D602D5",
x"02F402F302F202F102F002EF02EE02ED02EC02EB02EA02E902E802E702E602E5",
x"0000000000000000030002FF02FE02FD02FC02FB02FA02F902F802F702F602F5",
x"0310030F030E030D030C030B030A030903080307030603050304030303020301",
x"0320031F031E031D031C031B031A031903180317031603150314031303120311",
x"0330032F032E032D032C032B032A032903280327032603250324032303220321",
x"0340033F033E033D033C033B033A033903380337033603350334033303320331",
x"034C034B034A0349034803470346034503440343034203410000000000000000",
x"035C035B035A0359035803570356035503540353035203510350034F034E034D",
x"036C036B036A0369036803670366036503640363036203610360035F035E035D",
x"037C037B037A0379037803770376037503740373037203710370036F036E036D",
x"0388038703860385038403830382038100000000000000000380037F037E037D",
x"039803970396039503940393039203910390038F038E038D038C038B038A0389",
x"03A803A703A603A503A403A303A203A103A0039F039E039D039C039B039A0399",
x"03B803B703B603B503B403B303B203B103B003AF03AE03AD03AC03AB03AA03A9",
x"03C403C303C203C1000000000000000003C003BF03BE03BD03BC03BB03BA03B9",
x"03D403D303D203D103D003CF03CE03CD03CC03CB03CA03C903C803C703C603C5",
x"03E403E303E203E103E003DF03DE03DD03DC03DB03DA03D903D803D703D603D5",
x"03F403F303F203F103F003EF03EE03ED03EC03EB03EA03E903E803E703E603E5",
x"0000000000000000040003FF03FE03FD03FC03FB03FA03F903F803F703F603F5",
x"0410040F040E040D040C040B040A040904080407040604050404040304020401",
x"0420041F041E041D041C041B041A041904180417041604150414041304120411",
x"0430042F042E042D042C042B042A042904280427042604250424042304220421",
x"0440043F043E043D043C043B043A043904380437043604350434043304320431",
x"044C044B044A0449044804470446044504440443044204410000000000000000",
x"045C045B045A0459045804570456045504540453045204510450044F044E044D",
x"046C046B046A0469046804670466046504640463046204610460045F045E045D",
x"047C047B047A0479047804770476047504740473047204710470046F046E046D",
x"0488048704860485048404830482048100000000000000000480047F047E047D",
x"049804970496049504940493049204910490048F048E048D048C048B048A0489",
x"04A804A704A604A504A404A304A204A104A0049F049E049D049C049B049A0499",
x"04B804B704B604B504B404B304B204B104B004AF04AE04AD04AC04AB04AA04A9",
x"04C404C304C204C1FFFFFFFFFFFFFFFF04C004BF04BE04BD04BC04BB04BA04B9",
x"04D404D304D204D104D004CF04CE04CD04CC04CB04CA04C904C804C704C604C5",
x"0000000004E204E104E004DF04DE04DD04DC04DB04DA04D904D804D704D604D5",
x"0000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000"
	);                                  -- with data

begin

	p_comm_tb_avs_left_read_stimuli : process(clk_i, rst_i) is
		procedure p_readdata(read_address_i : std_logic_vector) is
			variable v_read_word_addr : natural range 0 to (c_CCD_IMGDATA_LENGTH - 1) := 0;
		begin

			-- set read word addr
			v_read_word_addr := to_integer(unsigned(read_address_i((g_ADDRESS_WIDTH - 1) downto 5))) mod (c_CCD_IMGDATA_LENGTH);

			-- check what imgdata selection is to be used
			if (c_CCD_IMGDATA_SELECTION = '0') then -- '0' = No Data / '1' = With Data
				-- imgdata selection is "No Data"
				-- return imgdata
				avs_avalon_mm_readata_o <= c_CCD_IMGDATA_NO_DATA(v_read_word_addr);
			else
				-- imgdata selection is "With Data"
				-- return imgdata
				avs_avalon_mm_readata_o <= c_CCD_IMGDATA_WITH_DATA(v_read_word_addr);
			end if;

		end procedure p_readdata;

	begin
		if (rst_i = '1') then
			avs_avalon_mm_readata_o     <= (others => '0');
			avs_avalon_mm_waitrequest_o <= '1';
		elsif (rising_edge(clk_i)) then
			avs_avalon_mm_readata_o     <= (others => '0');
			avs_avalon_mm_waitrequest_o <= '1';
			if (avs_avalon_mm_read_i = '1') then
				avs_avalon_mm_waitrequest_o <= '0';
				p_readdata(avs_avalon_mm_address_i);
			end if;
		end if;
	end process p_comm_tb_avs_left_read_stimuli;

end architecture RTL;
