-- MebX_Qsys_Project.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project is
	port (
		button_export                                                                           : in    std_logic_vector(3 downto 0)  := (others => '0'); --                                                       button.export
		clk50_clk                                                                               : in    std_logic                     := '0';             --                                                        clk50.clk
		comm_1_data_control_data_hold_signal                                                    : in    std_logic                     := '0';             --                                          comm_1_data_control.data_hold_signal
		comm_1_measurements_measurements_signal                                                 : out   std_logic_vector(7 downto 0);                     --                                          comm_1_measurements.measurements_signal
		comm_1_sync_sync_signal                                                                 : in    std_logic                     := '0';             --                                                  comm_1_sync.sync_signal
		comm_2_data_control_data_hold_signal                                                    : in    std_logic                     := '0';             --                                          comm_2_data_control.data_hold_signal
		comm_2_measurements_measurements_signal                                                 : out   std_logic_vector(7 downto 0);                     --                                          comm_2_measurements.measurements_signal
		comm_2_sync_sync_signal                                                                 : in    std_logic                     := '0';             --                                                  comm_2_sync.sync_signal
		comm_3_data_control_data_hold_signal                                                    : in    std_logic                     := '0';             --                                          comm_3_data_control.data_hold_signal
		comm_3_measurements_measurements_signal                                                 : out   std_logic_vector(7 downto 0);                     --                                          comm_3_measurements.measurements_signal
		comm_3_sync_sync_signal                                                                 : in    std_logic                     := '0';             --                                                  comm_3_sync.sync_signal
		comm_4_data_control_data_hold_signal                                                    : in    std_logic                     := '0';             --                                          comm_4_data_control.data_hold_signal
		comm_4_measurements_measurements_signal                                                 : out   std_logic_vector(7 downto 0);                     --                                          comm_4_measurements.measurements_signal
		comm_4_sync_sync_signal                                                                 : in    std_logic                     := '0';             --                                                  comm_4_sync.sync_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_echo_en_signal                    : out   std_logic;                                        --        communication_module_v2_ch1_conduit_end_rmap_echo_out.echo_en_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_echo_id_en_signal                 : out   std_logic;                                        --                                                             .echo_id_en_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrflag_signal             : out   std_logic;                                        --                                                             .in_fifo_wrflag_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrdata_signal             : out   std_logic_vector(7 downto 0);                     --                                                             .in_fifo_wrdata_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrreq_signal              : out   std_logic;                                        --                                                             .in_fifo_wrreq_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrflag_signal            : out   std_logic;                                        --                                                             .out_fifo_wrflag_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrdata_signal            : out   std_logic_vector(7 downto 0);                     --                                                             .out_fifo_wrdata_signal
		communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrreq_signal             : out   std_logic;                                        --                                                             .out_fifo_wrreq_signal
		communication_module_v2_ch2_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal : out   std_logic_vector(63 downto 0);                    -- communication_module_v2_ch2_conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_echo_en_signal                    : out   std_logic;                                        --        communication_module_v2_ch2_conduit_end_rmap_echo_out.echo_en_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_echo_id_en_signal                 : out   std_logic;                                        --                                                             .echo_id_en_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrflag_signal             : out   std_logic;                                        --                                                             .in_fifo_wrflag_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrdata_signal             : out   std_logic_vector(7 downto 0);                     --                                                             .in_fifo_wrdata_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrreq_signal              : out   std_logic;                                        --                                                             .in_fifo_wrreq_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrflag_signal            : out   std_logic;                                        --                                                             .out_fifo_wrflag_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrdata_signal            : out   std_logic_vector(7 downto 0);                     --                                                             .out_fifo_wrdata_signal
		communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrreq_signal             : out   std_logic;                                        --                                                             .out_fifo_wrreq_signal
		communication_module_v2_ch3_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal : out   std_logic_vector(63 downto 0);                    -- communication_module_v2_ch3_conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_echo_en_signal                    : out   std_logic;                                        --        communication_module_v2_ch3_conduit_end_rmap_echo_out.echo_en_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_echo_id_en_signal                 : out   std_logic;                                        --                                                             .echo_id_en_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrflag_signal             : out   std_logic;                                        --                                                             .in_fifo_wrflag_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrdata_signal             : out   std_logic_vector(7 downto 0);                     --                                                             .in_fifo_wrdata_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrreq_signal              : out   std_logic;                                        --                                                             .in_fifo_wrreq_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrflag_signal            : out   std_logic;                                        --                                                             .out_fifo_wrflag_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrdata_signal            : out   std_logic_vector(7 downto 0);                     --                                                             .out_fifo_wrdata_signal
		communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrreq_signal             : out   std_logic;                                        --                                                             .out_fifo_wrreq_signal
		communication_module_v2_ch4_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal : out   std_logic_vector(63 downto 0);                    -- communication_module_v2_ch4_conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_echo_en_signal                    : out   std_logic;                                        --        communication_module_v2_ch4_conduit_end_rmap_echo_out.echo_en_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_echo_id_en_signal                 : out   std_logic;                                        --                                                             .echo_id_en_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrflag_signal             : out   std_logic;                                        --                                                             .in_fifo_wrflag_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrdata_signal             : out   std_logic_vector(7 downto 0);                     --                                                             .in_fifo_wrdata_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrreq_signal              : out   std_logic;                                        --                                                             .in_fifo_wrreq_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrflag_signal            : out   std_logic;                                        --                                                             .out_fifo_wrflag_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrdata_signal            : out   std_logic_vector(7 downto 0);                     --                                                             .out_fifo_wrdata_signal
		communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrreq_signal             : out   std_logic;                                        --                                                             .out_fifo_wrreq_signal
		csense_adc_fo_export                                                                    : out   std_logic;                                        --                                                csense_adc_fo.export
		csense_cs_n_export                                                                      : out   std_logic_vector(1 downto 0);                     --                                                  csense_cs_n.export
		csense_sck_export                                                                       : out   std_logic;                                        --                                                   csense_sck.export
		csense_sdi_export                                                                       : out   std_logic;                                        --                                                   csense_sdi.export
		csense_sdo_export                                                                       : in    std_logic                     := '0';             --                                                   csense_sdo.export
		ctrl_io_lvds_export                                                                     : out   std_logic_vector(3 downto 0);                     --                                                 ctrl_io_lvds.export
		dip_export                                                                              : in    std_logic_vector(7 downto 0)  := (others => '0'); --                                                          dip.export
		ext_export                                                                              : in    std_logic                     := '0';             --                                                          ext.export
		ftdi_clk_clk                                                                            : in    std_logic                     := '0';             --                                                     ftdi_clk.clk
		ftdi_data_control_sync_pulse_signal                                                     : in    std_logic                     := '0';             --                                            ftdi_data_control.sync_pulse_signal
		ftdi_data_control_data_hold_signal                                                      : out   std_logic;                                        --                                                             .data_hold_signal
		led_de4_export                                                                          : out   std_logic_vector(7 downto 0);                     --                                                      led_de4.export
		led_painel_export                                                                       : out   std_logic_vector(20 downto 0);                    --                                                   led_painel.export
		m1_ddr2_i2c_scl_export                                                                  : out   std_logic;                                        --                                              m1_ddr2_i2c_scl.export
		m1_ddr2_i2c_sda_export                                                                  : inout std_logic                     := '0';             --                                              m1_ddr2_i2c_sda.export
		m1_ddr2_memory_mem_a                                                                    : out   std_logic_vector(13 downto 0);                    --                                               m1_ddr2_memory.mem_a
		m1_ddr2_memory_mem_ba                                                                   : out   std_logic_vector(2 downto 0);                     --                                                             .mem_ba
		m1_ddr2_memory_mem_ck                                                                   : out   std_logic_vector(1 downto 0);                     --                                                             .mem_ck
		m1_ddr2_memory_mem_ck_n                                                                 : out   std_logic_vector(1 downto 0);                     --                                                             .mem_ck_n
		m1_ddr2_memory_mem_cke                                                                  : out   std_logic_vector(1 downto 0);                     --                                                             .mem_cke
		m1_ddr2_memory_mem_cs_n                                                                 : out   std_logic_vector(1 downto 0);                     --                                                             .mem_cs_n
		m1_ddr2_memory_mem_dm                                                                   : out   std_logic_vector(7 downto 0);                     --                                                             .mem_dm
		m1_ddr2_memory_mem_ras_n                                                                : out   std_logic_vector(0 downto 0);                     --                                                             .mem_ras_n
		m1_ddr2_memory_mem_cas_n                                                                : out   std_logic_vector(0 downto 0);                     --                                                             .mem_cas_n
		m1_ddr2_memory_mem_we_n                                                                 : out   std_logic_vector(0 downto 0);                     --                                                             .mem_we_n
		m1_ddr2_memory_mem_dq                                                                   : inout std_logic_vector(63 downto 0) := (others => '0'); --                                                             .mem_dq
		m1_ddr2_memory_mem_dqs                                                                  : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                                             .mem_dqs
		m1_ddr2_memory_mem_dqs_n                                                                : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                                             .mem_dqs_n
		m1_ddr2_memory_mem_odt                                                                  : out   std_logic_vector(1 downto 0);                     --                                                             .mem_odt
		m1_ddr2_memory_pll_ref_clk_clk                                                          : in    std_logic                     := '0';             --                                   m1_ddr2_memory_pll_ref_clk.clk
		m1_ddr2_memory_status_local_init_done                                                   : out   std_logic;                                        --                                        m1_ddr2_memory_status.local_init_done
		m1_ddr2_memory_status_local_cal_success                                                 : out   std_logic;                                        --                                                             .local_cal_success
		m1_ddr2_memory_status_local_cal_fail                                                    : out   std_logic;                                        --                                                             .local_cal_fail
		m1_ddr2_oct_rdn                                                                         : in    std_logic                     := '0';             --                                                  m1_ddr2_oct.rdn
		m1_ddr2_oct_rup                                                                         : in    std_logic                     := '0';             --                                                             .rup
		m2_ddr2_i2c_scl_export                                                                  : out   std_logic;                                        --                                              m2_ddr2_i2c_scl.export
		m2_ddr2_i2c_sda_export                                                                  : inout std_logic                     := '0';             --                                              m2_ddr2_i2c_sda.export
		m2_ddr2_memory_mem_a                                                                    : out   std_logic_vector(13 downto 0);                    --                                               m2_ddr2_memory.mem_a
		m2_ddr2_memory_mem_ba                                                                   : out   std_logic_vector(2 downto 0);                     --                                                             .mem_ba
		m2_ddr2_memory_mem_ck                                                                   : out   std_logic_vector(1 downto 0);                     --                                                             .mem_ck
		m2_ddr2_memory_mem_ck_n                                                                 : out   std_logic_vector(1 downto 0);                     --                                                             .mem_ck_n
		m2_ddr2_memory_mem_cke                                                                  : out   std_logic_vector(1 downto 0);                     --                                                             .mem_cke
		m2_ddr2_memory_mem_cs_n                                                                 : out   std_logic_vector(1 downto 0);                     --                                                             .mem_cs_n
		m2_ddr2_memory_mem_dm                                                                   : out   std_logic_vector(7 downto 0);                     --                                                             .mem_dm
		m2_ddr2_memory_mem_ras_n                                                                : out   std_logic_vector(0 downto 0);                     --                                                             .mem_ras_n
		m2_ddr2_memory_mem_cas_n                                                                : out   std_logic_vector(0 downto 0);                     --                                                             .mem_cas_n
		m2_ddr2_memory_mem_we_n                                                                 : out   std_logic_vector(0 downto 0);                     --                                                             .mem_we_n
		m2_ddr2_memory_mem_dq                                                                   : inout std_logic_vector(63 downto 0) := (others => '0'); --                                                             .mem_dq
		m2_ddr2_memory_mem_dqs                                                                  : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                                             .mem_dqs
		m2_ddr2_memory_mem_dqs_n                                                                : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                                             .mem_dqs_n
		m2_ddr2_memory_mem_odt                                                                  : out   std_logic_vector(1 downto 0);                     --                                                             .mem_odt
		m2_ddr2_memory_dll_sharing_dll_pll_locked                                               : in    std_logic                     := '0';             --                                   m2_ddr2_memory_dll_sharing.dll_pll_locked
		m2_ddr2_memory_dll_sharing_dll_delayctrl                                                : out   std_logic_vector(5 downto 0);                     --                                                             .dll_delayctrl
		m2_ddr2_memory_pll_sharing_pll_mem_clk                                                  : out   std_logic;                                        --                                   m2_ddr2_memory_pll_sharing.pll_mem_clk
		m2_ddr2_memory_pll_sharing_pll_write_clk                                                : out   std_logic;                                        --                                                             .pll_write_clk
		m2_ddr2_memory_pll_sharing_pll_locked                                                   : out   std_logic;                                        --                                                             .pll_locked
		m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk                                    : out   std_logic;                                        --                                                             .pll_write_clk_pre_phy_clk
		m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk                                             : out   std_logic;                                        --                                                             .pll_addr_cmd_clk
		m2_ddr2_memory_pll_sharing_pll_avl_clk                                                  : out   std_logic;                                        --                                                             .pll_avl_clk
		m2_ddr2_memory_pll_sharing_pll_config_clk                                               : out   std_logic;                                        --                                                             .pll_config_clk
		m2_ddr2_memory_status_local_init_done                                                   : out   std_logic;                                        --                                        m2_ddr2_memory_status.local_init_done
		m2_ddr2_memory_status_local_cal_success                                                 : out   std_logic;                                        --                                                             .local_cal_success
		m2_ddr2_memory_status_local_cal_fail                                                    : out   std_logic;                                        --                                                             .local_cal_fail
		m2_ddr2_oct_rdn                                                                         : in    std_logic                     := '0';             --                                                  m2_ddr2_oct.rdn
		m2_ddr2_oct_rup                                                                         : in    std_logic                     := '0';             --                                                             .rup
		pio_ftdi_umft601a_module_reset_export                                                   : out   std_logic;                                        --                               pio_ftdi_umft601a_module_reset.export
		pio_iso_logic_signal_enable_export                                                      : out   std_logic;                                        --                                  pio_iso_logic_signal_enable.export
		pio_spw_demux_ch_1_select_export                                                        : out   std_logic_vector(1 downto 0);                     --                                    pio_spw_demux_ch_1_select.export
		pio_spw_demux_ch_2_select_export                                                        : out   std_logic_vector(1 downto 0);                     --                                    pio_spw_demux_ch_2_select.export
		pio_spw_demux_ch_3_select_export                                                        : out   std_logic_vector(1 downto 0);                     --                                    pio_spw_demux_ch_3_select.export
		pio_spw_demux_ch_4_select_export                                                        : out   std_logic_vector(1 downto 0);                     --                                    pio_spw_demux_ch_4_select.export
		rs232_uart_rxd                                                                          : in    std_logic                     := '0';             --                                                   rs232_uart.rxd
		rs232_uart_txd                                                                          : out   std_logic;                                        --                                                             .txd
		rst_reset_n                                                                             : in    std_logic                     := '0';             --                                                          rst.reset_n
		rst_controller_conduit_reset_input_t_reset_input_signal                                 : in    std_logic                     := '0';             --                           rst_controller_conduit_reset_input.t_reset_input_signal
		rst_controller_conduit_simucam_reset_t_simucam_reset_signal                             : out   std_logic;                                        --                         rst_controller_conduit_simucam_reset.t_simucam_reset_signal
		rtcc_alarm_export                                                                       : in    std_logic                     := '0';             --                                                   rtcc_alarm.export
		rtcc_cs_n_export                                                                        : out   std_logic;                                        --                                                    rtcc_cs_n.export
		rtcc_sck_export                                                                         : out   std_logic;                                        --                                                     rtcc_sck.export
		rtcc_sdi_export                                                                         : out   std_logic;                                        --                                                     rtcc_sdi.export
		rtcc_sdo_export                                                                         : in    std_logic                     := '0';             --                                                     rtcc_sdo.export
		sd_card_ip_b_SD_cmd                                                                     : inout std_logic                     := '0';             --                                                   sd_card_ip.b_SD_cmd
		sd_card_ip_b_SD_dat                                                                     : inout std_logic                     := '0';             --                                                             .b_SD_dat
		sd_card_ip_b_SD_dat3                                                                    : inout std_logic                     := '0';             --                                                             .b_SD_dat3
		sd_card_ip_o_SD_clock                                                                   : out   std_logic;                                        --                                                             .o_SD_clock
		sd_card_wp_n_io_export                                                                  : in    std_logic                     := '0';             --                                              sd_card_wp_n_io.export
		spwc_a_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_a_enable.spw_rx_enable_signal
		spwc_a_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_a_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_a_leds.spw_red_status_led_signal
		spwc_a_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_a_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_a_lvds.spw_lvds_p_data_in_signal
		spwc_a_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_a_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_a_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_a_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_a_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_a_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_a_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_b_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_b_enable.spw_rx_enable_signal
		spwc_b_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_b_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_b_leds.spw_red_status_led_signal
		spwc_b_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_b_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_b_lvds.spw_lvds_p_data_in_signal
		spwc_b_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_b_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_b_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_b_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_b_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_b_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_b_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_c_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_c_enable.spw_rx_enable_signal
		spwc_c_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_c_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_c_leds.spw_red_status_led_signal
		spwc_c_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_c_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_c_lvds.spw_lvds_p_data_in_signal
		spwc_c_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_c_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_c_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_c_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_c_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_c_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_c_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_d_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_d_enable.spw_rx_enable_signal
		spwc_d_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_d_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_d_leds.spw_red_status_led_signal
		spwc_d_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_d_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_d_lvds.spw_lvds_p_data_in_signal
		spwc_d_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_d_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_d_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_d_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_d_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_d_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_d_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_e_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_e_enable.spw_rx_enable_signal
		spwc_e_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_e_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_e_leds.spw_red_status_led_signal
		spwc_e_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_e_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_e_lvds.spw_lvds_p_data_in_signal
		spwc_e_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_e_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_e_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_e_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_e_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_e_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_e_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_f_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_f_enable.spw_rx_enable_signal
		spwc_f_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_f_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_f_leds.spw_red_status_led_signal
		spwc_f_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_f_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_f_lvds.spw_lvds_p_data_in_signal
		spwc_f_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_f_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_f_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_f_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_f_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_f_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_f_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_g_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_g_enable.spw_rx_enable_signal
		spwc_g_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_g_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_g_leds.spw_red_status_led_signal
		spwc_g_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_g_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_g_lvds.spw_lvds_p_data_in_signal
		spwc_g_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_g_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_g_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_g_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_g_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_g_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_g_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwc_h_enable_spw_rx_enable_signal                                                      : in    std_logic                     := '0';             --                                                spwc_h_enable.spw_rx_enable_signal
		spwc_h_enable_spw_tx_enable_signal                                                      : in    std_logic                     := '0';             --                                                             .spw_tx_enable_signal
		spwc_h_leds_spw_red_status_led_signal                                                   : out   std_logic;                                        --                                                  spwc_h_leds.spw_red_status_led_signal
		spwc_h_leds_spw_green_status_led_signal                                                 : out   std_logic;                                        --                                                             .spw_green_status_led_signal
		spwc_h_lvds_spw_lvds_p_data_in_signal                                                   : in    std_logic                     := '0';             --                                                  spwc_h_lvds.spw_lvds_p_data_in_signal
		spwc_h_lvds_spw_lvds_n_data_in_signal                                                   : in    std_logic                     := '0';             --                                                             .spw_lvds_n_data_in_signal
		spwc_h_lvds_spw_lvds_p_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_p_data_out_signal
		spwc_h_lvds_spw_lvds_n_data_out_signal                                                  : out   std_logic;                                        --                                                             .spw_lvds_n_data_out_signal
		spwc_h_lvds_spw_lvds_p_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_p_strobe_out_signal
		spwc_h_lvds_spw_lvds_n_strobe_out_signal                                                : out   std_logic;                                        --                                                             .spw_lvds_n_strobe_out_signal
		spwc_h_lvds_spw_lvds_p_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_p_strobe_in_signal
		spwc_h_lvds_spw_lvds_n_strobe_in_signal                                                 : in    std_logic                     := '0';             --                                                             .spw_lvds_n_strobe_in_signal
		spwd_ch1_select_demux_select_signal                                                     : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                              spwd_ch1_select.demux_select_signal
		spwd_ch2_select_demux_select_signal                                                     : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                              spwd_ch2_select.demux_select_signal
		spwd_ch3_select_demux_select_signal                                                     : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                              spwd_ch3_select.demux_select_signal
		spwd_ch4_select_demux_select_signal                                                     : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                              spwd_ch4_select.demux_select_signal
		sync_in_conduit                                                                         : in    std_logic                     := '0';             --                                                      sync_in.conduit
		sync_in_en_conduit                                                                      : in    std_logic                     := '0';             --                                                   sync_in_en.conduit
		sync_out_conduit                                                                        : out   std_logic;                                        --                                                     sync_out.conduit
		sync_out_en_conduit                                                                     : in    std_logic                     := '0';             --                                                  sync_out_en.conduit
		sync_spw1_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw1.conduit
		sync_spw2_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw2.conduit
		sync_spw3_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw3.conduit
		sync_spw4_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw4.conduit
		sync_spw5_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw5.conduit
		sync_spw6_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw6.conduit
		sync_spw7_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw7.conduit
		sync_spw8_conduit                                                                       : out   std_logic;                                        --                                                    sync_spw8.conduit
		temp_scl_export                                                                         : out   std_logic;                                        --                                                     temp_scl.export
		temp_sda_export                                                                         : inout std_logic                     := '0';             --                                                     temp_sda.export
		timer_1ms_external_port_export                                                          : out   std_logic;                                        --                                      timer_1ms_external_port.export
		timer_1us_external_port_export                                                          : out   std_logic;                                        --                                      timer_1us_external_port.export
		tristate_conduit_tcm_address_out                                                        : out   std_logic_vector(25 downto 0);                    --                                             tristate_conduit.tcm_address_out
		tristate_conduit_tcm_read_n_out                                                         : out   std_logic_vector(0 downto 0);                     --                                                             .tcm_read_n_out
		tristate_conduit_tcm_write_n_out                                                        : out   std_logic_vector(0 downto 0);                     --                                                             .tcm_write_n_out
		tristate_conduit_tcm_data_out                                                           : inout std_logic_vector(15 downto 0) := (others => '0'); --                                                             .tcm_data_out
		tristate_conduit_tcm_chipselect_n_out                                                   : out   std_logic_vector(0 downto 0);                     --                                                             .tcm_chipselect_n_out
		umft601a_pins_umft_clock_signal                                                         : in    std_logic                     := '0';             --                                                umft601a_pins.umft_clock_signal
		umft601a_pins_umft_txe_n_signal                                                         : in    std_logic                     := '0';             --                                                             .umft_txe_n_signal
		umft601a_pins_umft_rxf_n_signal                                                         : in    std_logic                     := '0';             --                                                             .umft_rxf_n_signal
		umft601a_pins_umft_data_signal                                                          : inout std_logic_vector(31 downto 0) := (others => '0'); --                                                             .umft_data_signal
		umft601a_pins_umft_be_signal                                                            : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                                             .umft_be_signal
		umft601a_pins_umft_wakeup_n_signal                                                      : inout std_logic                     := '0';             --                                                             .umft_wakeup_n_signal
		umft601a_pins_umft_gpio_bus_signal                                                      : inout std_logic_vector(1 downto 0)  := (others => '0'); --                                                             .umft_gpio_bus_signal
		umft601a_pins_umft_reset_n_signal                                                       : out   std_logic;                                        --                                                             .umft_reset_n_signal
		umft601a_pins_umft_wr_n_signal                                                          : out   std_logic;                                        --                                                             .umft_wr_n_signal
		umft601a_pins_umft_rd_n_signal                                                          : out   std_logic;                                        --                                                             .umft_rd_n_signal
		umft601a_pins_umft_oe_n_signal                                                          : out   std_logic;                                        --                                                             .umft_oe_n_signal
		umft601a_pins_umft_siwu_n_signal                                                        : out   std_logic                                         --                                                             .umft_siwu_n_signal
	);
end entity MebX_Qsys_Project;

architecture rtl of MebX_Qsys_Project is
	component Altera_UP_SD_Card_Avalon_Interface is
		port (
			i_avalon_chip_select : in    std_logic                     := 'X';             -- chipselect
			i_avalon_address     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			i_avalon_read        : in    std_logic                     := 'X';             -- read
			i_avalon_write       : in    std_logic                     := 'X';             -- write
			i_avalon_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest : out   std_logic;                                        -- waitrequest
			i_clock              : in    std_logic                     := 'X';             -- clk
			i_reset_n            : in    std_logic                     := 'X';             -- reset_n
			b_SD_cmd             : inout std_logic                     := 'X';             -- export
			b_SD_dat             : inout std_logic                     := 'X';             -- export
			b_SD_dat3            : inout std_logic                     := 'X';             -- export
			o_SD_clock           : out   std_logic                                         -- export
		);
	end component Altera_UP_SD_Card_Avalon_Interface;

	component comm_v2_top is
		port (
			reset_sink_reset_i                     : in  std_logic                      := 'X';             -- reset
			clock_sink_clk_i                       : in  std_logic                      := 'X';             -- clk
			channel_sync_i                         : in  std_logic                      := 'X';             -- sync_signal
			avs_config_address_i                   : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avs_config_write_i                     : in  std_logic                      := 'X';             -- write
			avs_config_writedata_i                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avs_config_read_i                      : in  std_logic                      := 'X';             -- read
			avs_config_readdata_o                  : out std_logic_vector(31 downto 0);                     -- readdata
			avs_config_waitrequest_o               : out std_logic;                                         -- waitrequest
			avm_left_buffer_readdata_i             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			avm_left_buffer_waitrequest_i          : in  std_logic                      := 'X';             -- waitrequest
			avm_left_buffer_address_o              : out std_logic_vector(63 downto 0);                     -- address
			avm_left_buffer_read_o                 : out std_logic;                                         -- read
			avm_right_buffer_readdata_i            : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			avm_right_buffer_waitrequest_i         : in  std_logic                      := 'X';             -- waitrequest
			avm_right_buffer_address_o             : out std_logic_vector(63 downto 0);                     -- address
			avm_right_buffer_read_o                : out std_logic;                                         -- read
			feeb_interrupt_sender_irq_o            : out std_logic;                                         -- irq
			rmap_interrupt_sender_irq_o            : out std_logic;                                         -- irq
			spw_link_status_started_i              : in  std_logic                      := 'X';             -- spw_link_status_started_signal
			spw_link_status_connecting_i           : in  std_logic                      := 'X';             -- spw_link_status_connecting_signal
			spw_link_status_running_i              : in  std_logic                      := 'X';             -- spw_link_status_running_signal
			spw_link_error_errdisc_i               : in  std_logic                      := 'X';             -- spw_link_error_errdisc_signal
			spw_link_error_errpar_i                : in  std_logic                      := 'X';             -- spw_link_error_errpar_signal
			spw_link_error_erresc_i                : in  std_logic                      := 'X';             -- spw_link_error_erresc_signal
			spw_link_error_errcred_i               : in  std_logic                      := 'X';             -- spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_i             : in  std_logic                      := 'X';             -- spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_i             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_i             : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_i           : in  std_logic                      := 'X';             -- spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_i           : in  std_logic                      := 'X';             -- spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_i            : in  std_logic                      := 'X';             -- spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_i            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_i             : in  std_logic                      := 'X';             -- spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_i           : in  std_logic                      := 'X';             -- spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_i          : in  std_logic                      := 'X';             -- spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_i         : in  std_logic                      := 'X';             -- spw_errinj_ctrl_errinj_ready_signal
			spw_link_command_enable_o              : out std_logic;                                         -- spw_link_command_enable_signal
			spw_link_command_autostart_o           : out std_logic;                                         -- spw_link_command_autostart_signal
			spw_link_command_linkstart_o           : out std_logic;                                         -- spw_link_command_linkstart_signal
			spw_link_command_linkdis_o             : out std_logic;                                         -- spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_o            : out std_logic_vector(7 downto 0);                      -- spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_o              : out std_logic;                                         -- spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_o              : out std_logic_vector(1 downto 0);                      -- spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_o              : out std_logic_vector(5 downto 0);                      -- spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_o           : out std_logic;                                         -- spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_o          : out std_logic;                                         -- spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_o           : out std_logic;                                         -- spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_o           : out std_logic_vector(7 downto 0);                      -- spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_o         : out std_logic;                                         -- spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_o         : out std_logic;                                         -- spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_o          : out std_logic_vector(3 downto 0);                      -- spw_errinj_ctrl_errinj_code_signal
			rmap_echo_echo_en_o                    : out std_logic;                                         -- echo_en_signal
			rmap_echo_echo_id_en_o                 : out std_logic;                                         -- echo_id_en_signal
			rmap_echo_in_fifo_wrflag_o             : out std_logic;                                         -- in_fifo_wrflag_signal
			rmap_echo_in_fifo_wrdata_o             : out std_logic_vector(7 downto 0);                      -- in_fifo_wrdata_signal
			rmap_echo_in_fifo_wrreq_o              : out std_logic;                                         -- in_fifo_wrreq_signal
			rmap_echo_out_fifo_wrflag_o            : out std_logic;                                         -- out_fifo_wrflag_signal
			rmap_echo_out_fifo_wrdata_o            : out std_logic_vector(7 downto 0);                      -- out_fifo_wrdata_signal
			rmap_echo_out_fifo_wrreq_o             : out std_logic;                                         -- out_fifo_wrreq_signal
			rmm_deb_rmap_target_wr_waitrequest_i   : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_deb_rmap_target_readdata_i         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_deb_rmap_target_rd_waitrequest_i   : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_deb_rmap_target_wr_address_o       : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_deb_rmap_target_write_o            : out std_logic;                                         -- write_signal
			rmm_deb_rmap_target_writedata_o        : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_deb_rmap_target_rd_address_o       : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_deb_rmap_target_read_o             : out std_logic;                                         -- read_signal
			rmm_deb_fee_hk_wr_waitrequest_i        : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_deb_fee_hk_readdata_i              : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_deb_fee_hk_rd_waitrequest_i        : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_deb_fee_hk_wr_address_o            : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_deb_fee_hk_write_o                 : out std_logic;                                         -- write_signal
			rmm_deb_fee_hk_writedata_o             : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_deb_fee_hk_rd_address_o            : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_deb_fee_hk_read_o                  : out std_logic;                                         -- read_signal
			rmm_aeb1_rmap_target_wr_waitrequest_i  : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb1_rmap_target_readdata_i        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb1_rmap_target_rd_waitrequest_i  : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb1_rmap_target_wr_address_o      : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb1_rmap_target_write_o           : out std_logic;                                         -- write_signal
			rmm_aeb1_rmap_target_writedata_o       : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb1_rmap_target_rd_address_o      : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb1_rmap_target_read_o            : out std_logic;                                         -- read_signal
			rmm_aeb1_fee_hk_wr_waitrequest_i       : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb1_fee_hk_readdata_i             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb1_fee_hk_rd_waitrequest_i       : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb1_fee_hk_wr_address_o           : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb1_fee_hk_write_o                : out std_logic;                                         -- write_signal
			rmm_aeb1_fee_hk_writedata_o            : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb1_fee_hk_rd_address_o           : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb1_fee_hk_read_o                 : out std_logic;                                         -- read_signal
			rmm_aeb2_rmap_target_wr_waitrequest_i  : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb2_rmap_target_readdata_i        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb2_rmap_target_rd_waitrequest_i  : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb2_rmap_target_wr_address_o      : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb2_rmap_target_write_o           : out std_logic;                                         -- write_signal
			rmm_aeb2_rmap_target_writedata_o       : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb2_rmap_target_rd_address_o      : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb2_rmap_target_read_o            : out std_logic;                                         -- read_signal
			rmm_aeb2_fee_hk_wr_waitrequest_i       : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb2_fee_hk_readdata_i             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb2_fee_hk_rd_waitrequest_i       : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb2_fee_hk_wr_address_o           : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb2_fee_hk_write_o                : out std_logic;                                         -- write_signal
			rmm_aeb2_fee_hk_writedata_o            : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb2_fee_hk_rd_address_o           : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb2_fee_hk_read_o                 : out std_logic;                                         -- read_signal
			rmm_aeb3_rmap_target_wr_waitrequest_i  : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb3_rmap_target_readdata_i        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb3_rmap_target_rd_waitrequest_i  : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb3_rmap_target_wr_address_o      : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb3_rmap_target_write_o           : out std_logic;                                         -- write_signal
			rmm_aeb3_rmap_target_writedata_o       : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb3_rmap_target_rd_address_o      : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb3_rmap_target_read_o            : out std_logic;                                         -- read_signal
			rmm_aeb3_fee_hk_wr_waitrequest_i       : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb3_fee_hk_readdata_i             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb3_fee_hk_rd_waitrequest_i       : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb3_fee_hk_wr_address_o           : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb3_fee_hk_write_o                : out std_logic;                                         -- write_signal
			rmm_aeb3_fee_hk_writedata_o            : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb3_fee_hk_rd_address_o           : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb3_fee_hk_read_o                 : out std_logic;                                         -- read_signal
			rmm_aeb4_rmap_target_wr_waitrequest_i  : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb4_rmap_target_readdata_i        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb4_rmap_target_rd_waitrequest_i  : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb4_rmap_target_wr_address_o      : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb4_rmap_target_write_o           : out std_logic;                                         -- write_signal
			rmm_aeb4_rmap_target_writedata_o       : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb4_rmap_target_rd_address_o      : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb4_rmap_target_read_o            : out std_logic;                                         -- read_signal
			rmm_aeb4_fee_hk_wr_waitrequest_i       : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			rmm_aeb4_fee_hk_readdata_i             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			rmm_aeb4_fee_hk_rd_waitrequest_i       : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			rmm_aeb4_fee_hk_wr_address_o           : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			rmm_aeb4_fee_hk_write_o                : out std_logic;                                         -- write_signal
			rmm_aeb4_fee_hk_writedata_o            : out std_logic_vector(7 downto 0);                      -- writedata_signal
			rmm_aeb4_fee_hk_rd_address_o           : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			rmm_aeb4_fee_hk_read_o                 : out std_logic;                                         -- read_signal
			channel_hk_rmap_target_status_o        : out std_logic_vector(7 downto 0);                      -- rmap_target_status_signal
			channel_hk_rmap_target_indicate_o      : out std_logic;                                         -- rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o       : out std_logic;                                         -- spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o       : out std_logic;                                         -- spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o       : out std_logic;                                         -- spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o       : out std_logic;                                         -- spw_link_disconnect_signal
			channel_hk_spw_link_started_o          : out std_logic;                                         -- spw_link_started_signal
			channel_hk_spw_link_connecting_o       : out std_logic;                                         -- spw_link_connecting_signal
			channel_hk_spw_link_running_o          : out std_logic;                                         -- spw_link_running_signal
			channel_hk_frame_counter_o             : out std_logic_vector(15 downto 0);                     -- frame_counter_signal
			channel_hk_left_buffer_ccd_number_o    : out std_logic_vector(1 downto 0);                      -- left_buffer_ccd_number_signal
			channel_hk_right_buffer_ccd_number_o   : out std_logic_vector(1 downto 0);                      -- right_buffer_ccd_number_signal
			channel_hk_left_buffer_ccd_side_o      : out std_logic;                                         -- left_buffer_ccd_side_signal
			channel_hk_right_buffer_ccd_side_o     : out std_logic;                                         -- right_buffer_ccd_side_signal
			channel_hk_err_left_buffer_overflow_o  : out std_logic;                                         -- err_left_buffer_overflow_signal
			channel_hk_err_right_buffer_overflow_o : out std_logic;                                         -- err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_o          : out std_logic_vector(63 downto 0);                     -- win_mem_addr_offset_signal
			comm_data_control_data_hold_i          : in  std_logic                      := 'X';             -- data_hold_signal
			comm_measurements_o                    : out std_logic_vector(7 downto 0)                       -- measurements_signal
		);
	end component comm_v2_top;

	component ftdi_usb3_top is
		port (
			clock_sink_clk_i                      : in    std_logic                      := 'X';             -- clk
			reset_sink_reset_i                    : in    std_logic                      := 'X';             -- reset
			umft601a_clock_sink_clk_i             : in    std_logic                      := 'X';             -- clk
			umft601a_clock_pin_i                  : in    std_logic                      := 'X';             -- umft_clock_signal
			umft601a_txe_n_pin_i                  : in    std_logic                      := 'X';             -- umft_txe_n_signal
			umft601a_rxf_n_pin_i                  : in    std_logic                      := 'X';             -- umft_rxf_n_signal
			umft601a_data_bus_io                  : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- umft_data_signal
			umft601a_be_bus_io                    : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- umft_be_signal
			umft601a_wakeup_n_pin_io              : inout std_logic                      := 'X';             -- umft_wakeup_n_signal
			umft601a_gpio_bus_io                  : inout std_logic_vector(1 downto 0)   := (others => 'X'); -- umft_gpio_bus_signal
			umft601a_reset_n_pin_o                : out   std_logic;                                         -- umft_reset_n_signal
			umft601a_wr_n_pin_o                   : out   std_logic;                                         -- umft_wr_n_signal
			umft601a_rd_n_pin_o                   : out   std_logic;                                         -- umft_rd_n_signal
			umft601a_oe_n_pin_o                   : out   std_logic;                                         -- umft_oe_n_signal
			umft601a_siwu_n_pin_o                 : out   std_logic;                                         -- umft_siwu_n_signal
			avalon_slave_config_address_i         : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avalon_slave_config_write_i           : in    std_logic                      := 'X';             -- write
			avalon_slave_config_writedata_i       : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avalon_slave_config_read_i            : in    std_logic                      := 'X';             -- read
			avalon_slave_config_readdata_o        : out   std_logic_vector(31 downto 0);                     -- readdata
			avalon_slave_config_waitrequest_o     : out   std_logic;                                         -- waitrequest
			avalon_master_data_readdata_i         : in    std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			avalon_master_data_waitrequest_i      : in    std_logic                      := 'X';             -- waitrequest
			avalon_master_data_address_o          : out   std_logic_vector(63 downto 0);                     -- address
			avalon_master_data_read_o             : out   std_logic;                                         -- read
			avalon_master_data_write_o            : out   std_logic;                                         -- write
			avalon_master_data_writedata_o        : out   std_logic_vector(255 downto 0);                    -- writedata
			avalon_imgt_master_data_waitrequest_i : in    std_logic                      := 'X';             -- waitrequest
			avalon_imgt_master_data_address_o     : out   std_logic_vector(63 downto 0);                     -- address
			avalon_imgt_master_data_write_o       : out   std_logic;                                         -- write
			avalon_imgt_master_data_writedata_o   : out   std_logic_vector(15 downto 0);                     -- writedata
			rx_interrupt_sender_irq_o             : out   std_logic;                                         -- irq
			tx_interrupt_sender_irq_o             : out   std_logic;                                         -- irq
			ftdi_data_control_sync_pulse_i        : in    std_logic                      := 'X';             -- sync_pulse_signal
			ftdi_data_control_data_hold_o         : out   std_logic                                          -- data_hold_signal
		);
	end component ftdi_usb3_top;

	component mfil_memory_filler_top is
		port (
			clock_sink_clk_i                  : in  std_logic                      := 'X';             -- clk
			reset_sink_reset_i                : in  std_logic                      := 'X';             -- reset
			avalon_slave_config_address_i     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avalon_slave_config_byteenable_i  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			avalon_slave_config_write_i       : in  std_logic                      := 'X';             -- write
			avalon_slave_config_writedata_i   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avalon_slave_config_read_i        : in  std_logic                      := 'X';             -- read
			avalon_slave_config_readdata_o    : out std_logic_vector(31 downto 0);                     -- readdata
			avalon_slave_config_waitrequest_o : out std_logic;                                         -- waitrequest
			avalon_master_data_waitrequest_i  : in  std_logic                      := 'X';             -- waitrequest
			avalon_master_data_address_o      : out std_logic_vector(63 downto 0);                     -- address
			avalon_master_data_write_o        : out std_logic;                                         -- write
			avalon_master_data_writedata_o    : out std_logic_vector(255 downto 0)                     -- writedata
		);
	end component mfil_memory_filler_top;

	component spwc_spacewire_channel_top is
		port (
			reset_i                        : in  std_logic                    := 'X';             -- reset
			clk_100_i                      : in  std_logic                    := 'X';             -- clk
			clk_200_i                      : in  std_logic                    := 'X';             -- clk
			spw_lvds_p_data_in_i           : in  std_logic                    := 'X';             -- spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           : in  std_logic                    := 'X';             -- spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          : out std_logic;                                       -- spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          : out std_logic;                                       -- spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        : out std_logic;                                       -- spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        : out std_logic;                                       -- spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         : in  std_logic                    := 'X';             -- spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         : in  std_logic                    := 'X';             -- spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                : in  std_logic                    := 'X';             -- spw_rx_enable_signal
			spw_tx_enable_i                : in  std_logic                    := 'X';             -- spw_tx_enable_signal
			spw_red_status_led_o           : out std_logic;                                       -- spw_red_status_led_signal
			spw_green_status_led_o         : out std_logic;                                       -- spw_green_status_led_signal
			spw_link_command_enable_i      : in  std_logic                    := 'X';             -- spw_link_command_enable_signal
			spw_link_command_autostart_i   : in  std_logic                    := 'X';             -- spw_link_command_autostart_signal
			spw_link_command_linkstart_i   : in  std_logic                    := 'X';             -- spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     : in  std_logic                    := 'X';             -- spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      : in  std_logic                    := 'X';             -- spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      : in  std_logic_vector(1 downto 0) := (others => 'X'); -- spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      : in  std_logic_vector(5 downto 0) := (others => 'X'); -- spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   : in  std_logic                    := 'X';             -- spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  : in  std_logic                    := 'X';             -- spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   : in  std_logic                    := 'X';             -- spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i : in  std_logic                    := 'X';             -- spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i : in  std_logic                    := 'X';             -- spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  : in  std_logic_vector(3 downto 0) := (others => 'X'); -- spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      : out std_logic;                                       -- spw_link_status_started_signal
			spw_link_status_connecting_o   : out std_logic;                                       -- spw_link_status_connecting_signal
			spw_link_status_running_o      : out std_logic;                                       -- spw_link_status_running_signal
			spw_link_error_errdisc_o       : out std_logic;                                       -- spw_link_error_errdisc_signal
			spw_link_error_errpar_o        : out std_logic;                                       -- spw_link_error_errpar_signal
			spw_link_error_erresc_o        : out std_logic;                                       -- spw_link_error_erresc_signal
			spw_link_error_errcred_o       : out std_logic;                                       -- spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     : out std_logic;                                       -- spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     : out std_logic_vector(1 downto 0);                    -- spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     : out std_logic_vector(5 downto 0);                    -- spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   : out std_logic;                                       -- spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   : out std_logic;                                       -- spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    : out std_logic;                                       -- spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    : out std_logic_vector(7 downto 0);                    -- spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     : out std_logic;                                       -- spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   : out std_logic;                                       -- spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  : out std_logic;                                       -- spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o : out std_logic                                        -- spw_errinj_ctrl_errinj_ready_signal
		);
	end component spwc_spacewire_channel_top;

	component spwd_spacewire_demux_top is
		port (
			reset_i                            : in  std_logic                    := 'X';             -- reset
			clock_i                            : in  std_logic                    := 'X';             -- clk
			demux_select_i                     : in  std_logic_vector(1 downto 0) := (others => 'X'); -- demux_select_signal
			spw_link_command_enable_i          : in  std_logic                    := 'X';             -- spw_link_command_enable_signal
			spw_link_command_autostart_i       : in  std_logic                    := 'X';             -- spw_link_command_autostart_signal
			spw_link_command_linkstart_i       : in  std_logic                    := 'X';             -- spw_link_command_linkstart_signal
			spw_link_command_linkdis_i         : in  std_logic                    := 'X';             -- spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i        : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i          : in  std_logic                    := 'X';             -- spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i          : in  std_logic_vector(1 downto 0) := (others => 'X'); -- spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i          : in  std_logic_vector(5 downto 0) := (others => 'X'); -- spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i       : in  std_logic                    := 'X';             -- spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i      : in  std_logic                    := 'X';             -- spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i       : in  std_logic                    := 'X';             -- spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i       : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i     : in  std_logic                    := 'X';             -- spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i     : in  std_logic                    := 'X';             -- spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i      : in  std_logic_vector(3 downto 0) := (others => 'X'); -- spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o          : out std_logic;                                       -- spw_link_status_started_signal
			spw_link_status_connecting_o       : out std_logic;                                       -- spw_link_status_connecting_signal
			spw_link_status_running_o          : out std_logic;                                       -- spw_link_status_running_signal
			spw_link_error_errdisc_o           : out std_logic;                                       -- spw_link_error_errdisc_signal
			spw_link_error_errpar_o            : out std_logic;                                       -- spw_link_error_errpar_signal
			spw_link_error_erresc_o            : out std_logic;                                       -- spw_link_error_erresc_signal
			spw_link_error_errcred_o           : out std_logic;                                       -- spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o         : out std_logic;                                       -- spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o         : out std_logic_vector(1 downto 0);                    -- spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o         : out std_logic_vector(5 downto 0);                    -- spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o       : out std_logic;                                       -- spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o       : out std_logic;                                       -- spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o        : out std_logic;                                       -- spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o        : out std_logic_vector(7 downto 0);                    -- spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o         : out std_logic;                                       -- spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o       : out std_logic;                                       -- spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o      : out std_logic;                                       -- spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o     : out std_logic;                                       -- spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_status_started_i      : in  std_logic                    := 'X';             -- spw_link_status_started_signal
			spw_ct0_link_status_connecting_i   : in  std_logic                    := 'X';             -- spw_link_status_connecting_signal
			spw_ct0_link_status_running_i      : in  std_logic                    := 'X';             -- spw_link_status_running_signal
			spw_ct0_link_error_errdisc_i       : in  std_logic                    := 'X';             -- spw_link_error_errdisc_signal
			spw_ct0_link_error_errpar_i        : in  std_logic                    := 'X';             -- spw_link_error_errpar_signal
			spw_ct0_link_error_erresc_i        : in  std_logic                    := 'X';             -- spw_link_error_erresc_signal
			spw_ct0_link_error_errcred_i       : in  std_logic                    := 'X';             -- spw_link_error_errcred_signal
			spw_ct0_timecode_rx_tick_out_i     : in  std_logic                    := 'X';             -- spw_timecode_rx_tick_out_signal
			spw_ct0_timecode_rx_ctrl_out_i     : in  std_logic_vector(1 downto 0) := (others => 'X'); -- spw_timecode_rx_ctrl_out_signal
			spw_ct0_timecode_rx_time_out_i     : in  std_logic_vector(5 downto 0) := (others => 'X'); -- spw_timecode_rx_time_out_signal
			spw_ct0_data_rx_status_rxvalid_i   : in  std_logic                    := 'X';             -- spw_data_rx_status_rxvalid_signal
			spw_ct0_data_rx_status_rxhalff_i   : in  std_logic                    := 'X';             -- spw_data_rx_status_rxhalff_signal
			spw_ct0_data_rx_status_rxflag_i    : in  std_logic                    := 'X';             -- spw_data_rx_status_rxflag_signal
			spw_ct0_data_rx_status_rxdata_i    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_data_rx_status_rxdata_signal
			spw_ct0_data_tx_status_txrdy_i     : in  std_logic                    := 'X';             -- spw_data_tx_status_txrdy_signal
			spw_ct0_data_tx_status_txhalff_i   : in  std_logic                    := 'X';             -- spw_data_tx_status_txhalff_signal
			spw_ct0_errinj_ctrl_errinj_busy_i  : in  std_logic                    := 'X';             -- spw_errinj_ctrl_errinj_busy_signal
			spw_ct0_errinj_ctrl_errinj_ready_i : in  std_logic                    := 'X';             -- spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_command_enable_o      : out std_logic;                                       -- spw_link_command_enable_signal
			spw_ct0_link_command_autostart_o   : out std_logic;                                       -- spw_link_command_autostart_signal
			spw_ct0_link_command_linkstart_o   : out std_logic;                                       -- spw_link_command_linkstart_signal
			spw_ct0_link_command_linkdis_o     : out std_logic;                                       -- spw_link_command_linkdis_signal
			spw_ct0_link_command_txdivcnt_o    : out std_logic_vector(7 downto 0);                    -- spw_link_command_txdivcnt_signal
			spw_ct0_timecode_tx_tick_in_o      : out std_logic;                                       -- spw_timecode_tx_tick_in_signal
			spw_ct0_timecode_tx_ctrl_in_o      : out std_logic_vector(1 downto 0);                    -- spw_timecode_tx_ctrl_in_signal
			spw_ct0_timecode_tx_time_in_o      : out std_logic_vector(5 downto 0);                    -- spw_timecode_tx_time_in_signal
			spw_ct0_data_rx_command_rxread_o   : out std_logic;                                       -- spw_data_rx_command_rxread_signal
			spw_ct0_data_tx_command_txwrite_o  : out std_logic;                                       -- spw_data_tx_command_txwrite_signal
			spw_ct0_data_tx_command_txflag_o   : out std_logic;                                       -- spw_data_tx_command_txflag_signal
			spw_ct0_data_tx_command_txdata_o   : out std_logic_vector(7 downto 0);                    -- spw_data_tx_command_txdata_signal
			spw_ct0_errinj_ctrl_start_errinj_o : out std_logic;                                       -- spw_errinj_ctrl_start_errinj_signal
			spw_ct0_errinj_ctrl_reset_errinj_o : out std_logic;                                       -- spw_errinj_ctrl_reset_errinj_signal
			spw_ct0_errinj_ctrl_errinj_code_o  : out std_logic_vector(3 downto 0);                    -- spw_errinj_ctrl_errinj_code_signal
			spw_ct1_link_status_started_i      : in  std_logic                    := 'X';             -- spw_link_status_started_signal
			spw_ct1_link_status_connecting_i   : in  std_logic                    := 'X';             -- spw_link_status_connecting_signal
			spw_ct1_link_status_running_i      : in  std_logic                    := 'X';             -- spw_link_status_running_signal
			spw_ct1_link_error_errdisc_i       : in  std_logic                    := 'X';             -- spw_link_error_errdisc_signal
			spw_ct1_link_error_errpar_i        : in  std_logic                    := 'X';             -- spw_link_error_errpar_signal
			spw_ct1_link_error_erresc_i        : in  std_logic                    := 'X';             -- spw_link_error_erresc_signal
			spw_ct1_link_error_errcred_i       : in  std_logic                    := 'X';             -- spw_link_error_errcred_signal
			spw_ct1_timecode_rx_tick_out_i     : in  std_logic                    := 'X';             -- spw_timecode_rx_tick_out_signal
			spw_ct1_timecode_rx_ctrl_out_i     : in  std_logic_vector(1 downto 0) := (others => 'X'); -- spw_timecode_rx_ctrl_out_signal
			spw_ct1_timecode_rx_time_out_i     : in  std_logic_vector(5 downto 0) := (others => 'X'); -- spw_timecode_rx_time_out_signal
			spw_ct1_data_rx_status_rxvalid_i   : in  std_logic                    := 'X';             -- spw_data_rx_status_rxvalid_signal
			spw_ct1_data_rx_status_rxhalff_i   : in  std_logic                    := 'X';             -- spw_data_rx_status_rxhalff_signal
			spw_ct1_data_rx_status_rxflag_i    : in  std_logic                    := 'X';             -- spw_data_rx_status_rxflag_signal
			spw_ct1_data_rx_status_rxdata_i    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- spw_data_rx_status_rxdata_signal
			spw_ct1_data_tx_status_txrdy_i     : in  std_logic                    := 'X';             -- spw_data_tx_status_txrdy_signal
			spw_ct1_data_tx_status_txhalff_i   : in  std_logic                    := 'X';             -- spw_data_tx_status_txhalff_signal
			spw_ct1_errinj_ctrl_errinj_busy_i  : in  std_logic                    := 'X';             -- spw_errinj_ctrl_errinj_busy_signal
			spw_ct1_errinj_ctrl_errinj_ready_i : in  std_logic                    := 'X';             -- spw_errinj_ctrl_errinj_ready_signal
			spw_ct1_link_command_enable_o      : out std_logic;                                       -- spw_link_command_enable_signal
			spw_ct1_link_command_autostart_o   : out std_logic;                                       -- spw_link_command_autostart_signal
			spw_ct1_link_command_linkstart_o   : out std_logic;                                       -- spw_link_command_linkstart_signal
			spw_ct1_link_command_linkdis_o     : out std_logic;                                       -- spw_link_command_linkdis_signal
			spw_ct1_link_command_txdivcnt_o    : out std_logic_vector(7 downto 0);                    -- spw_link_command_txdivcnt_signal
			spw_ct1_timecode_tx_tick_in_o      : out std_logic;                                       -- spw_timecode_tx_tick_in_signal
			spw_ct1_timecode_tx_ctrl_in_o      : out std_logic_vector(1 downto 0);                    -- spw_timecode_tx_ctrl_in_signal
			spw_ct1_timecode_tx_time_in_o      : out std_logic_vector(5 downto 0);                    -- spw_timecode_tx_time_in_signal
			spw_ct1_data_rx_command_rxread_o   : out std_logic;                                       -- spw_data_rx_command_rxread_signal
			spw_ct1_data_tx_command_txwrite_o  : out std_logic;                                       -- spw_data_tx_command_txwrite_signal
			spw_ct1_data_tx_command_txflag_o   : out std_logic;                                       -- spw_data_tx_command_txflag_signal
			spw_ct1_data_tx_command_txdata_o   : out std_logic_vector(7 downto 0);                    -- spw_data_tx_command_txdata_signal
			spw_ct1_errinj_ctrl_start_errinj_o : out std_logic;                                       -- spw_errinj_ctrl_start_errinj_signal
			spw_ct1_errinj_ctrl_reset_errinj_o : out std_logic;                                       -- spw_errinj_ctrl_reset_errinj_signal
			spw_ct1_errinj_ctrl_errinj_code_o  : out std_logic_vector(3 downto 0)                     -- spw_errinj_ctrl_errinj_code_signal
		);
	end component spwd_spacewire_demux_top;

	component MebX_Qsys_Project_csense_adc_fo is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_csense_adc_fo;

	component MebX_Qsys_Project_csense_cs_n is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_csense_cs_n;

	component MebX_Qsys_Project_csense_sdo is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_csense_sdo;

	component altera_address_span_extender is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			avs_s0_address       : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                     := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                     := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_readdatavalid : out std_logic;                                        -- readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_burstcount    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_m0_read          : out std_logic;                                        -- read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                        -- write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_m0_burstcount    : out std_logic_vector(7 downto 0);                     -- burstcount
			avs_cntl_read        : in  std_logic                     := 'X';             -- read
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);                    -- readdata
			avs_cntl_write       : in  std_logic                     := 'X';             -- write
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- address
		);
	end component altera_address_span_extender;

	component MebX_Qsys_Project_ext_flash is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(25 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component MebX_Qsys_Project_ext_flash;

	component MebX_Qsys_Project_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_jtag_uart_0;

	component MebX_Qsys_Project_m1_ddr2_i2c_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_m1_ddr2_i2c_sda;

	component MebX_Qsys_Project_m1_ddr2_memory is
		port (
			pll_ref_clk        : in    std_logic                      := 'X';             -- clk
			global_reset_n     : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n       : in    std_logic                      := 'X';             -- reset_n
			afi_clk            : out   std_logic;                                         -- clk
			afi_half_clk       : out   std_logic;                                         -- clk
			afi_reset_n        : out   std_logic;                                         -- reset_n
			afi_reset_export_n : out   std_logic;                                         -- reset_n
			mem_a              : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba             : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck             : out   std_logic_vector(1 downto 0);                      -- mem_ck
			mem_ck_n           : out   std_logic_vector(1 downto 0);                      -- mem_ck_n
			mem_cke            : out   std_logic_vector(1 downto 0);                      -- mem_cke
			mem_cs_n           : out   std_logic_vector(1 downto 0);                      -- mem_cs_n
			mem_dm             : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n          : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n          : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n           : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_dq             : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs            : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n          : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt            : out   std_logic_vector(1 downto 0);                      -- mem_odt
			avl_ready          : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin     : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr           : in    std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid    : out   std_logic;                                         -- readdatavalid
			avl_rdata          : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata          : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req       : in    std_logic                      := 'X';             -- read
			avl_write_req      : in    std_logic                      := 'X';             -- write
			avl_size           : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			local_init_done    : out   std_logic;                                         -- local_init_done
			local_cal_success  : out   std_logic;                                         -- local_cal_success
			local_cal_fail     : out   std_logic;                                         -- local_cal_fail
			oct_rdn            : in    std_logic                      := 'X';             -- rdn
			oct_rup            : in    std_logic                      := 'X'              -- rup
		);
	end component MebX_Qsys_Project_m1_ddr2_memory;

	component MebX_Qsys_Project_m2_ddr2_memory is
		port (
			pll_ref_clk               : in    std_logic                      := 'X';             -- clk
			global_reset_n            : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n              : in    std_logic                      := 'X';             -- reset_n
			afi_clk                   : out   std_logic;                                         -- clk
			afi_half_clk              : out   std_logic;                                         -- clk
			afi_reset_n               : out   std_logic;                                         -- reset_n
			afi_reset_export_n        : out   std_logic;                                         -- reset_n
			mem_a                     : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba                    : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                    : out   std_logic_vector(1 downto 0);                      -- mem_ck
			mem_ck_n                  : out   std_logic_vector(1 downto 0);                      -- mem_ck_n
			mem_cke                   : out   std_logic_vector(1 downto 0);                      -- mem_cke
			mem_cs_n                  : out   std_logic_vector(1 downto 0);                      -- mem_cs_n
			mem_dm                    : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n                 : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n                 : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n                  : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_dq                    : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                   : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                 : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                   : out   std_logic_vector(1 downto 0);                      -- mem_odt
			avl_ready                 : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin            : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr                  : in    std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid           : out   std_logic;                                         -- readdatavalid
			avl_rdata                 : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata                 : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be                    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req              : in    std_logic                      := 'X';             -- read
			avl_write_req             : in    std_logic                      := 'X';             -- write
			avl_size                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			local_init_done           : out   std_logic;                                         -- local_init_done
			local_cal_success         : out   std_logic;                                         -- local_cal_success
			local_cal_fail            : out   std_logic;                                         -- local_cal_fail
			oct_rdn                   : in    std_logic                      := 'X';             -- rdn
			oct_rup                   : in    std_logic                      := 'X';             -- rup
			pll_mem_clk               : out   std_logic;                                         -- pll_mem_clk
			pll_write_clk             : out   std_logic;                                         -- pll_write_clk
			pll_locked                : out   std_logic;                                         -- pll_locked
			pll_write_clk_pre_phy_clk : out   std_logic;                                         -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          : out   std_logic;                                         -- pll_addr_cmd_clk
			pll_avl_clk               : out   std_logic;                                         -- pll_avl_clk
			pll_config_clk            : out   std_logic;                                         -- pll_config_clk
			dll_pll_locked            : in    std_logic                      := 'X';             -- dll_pll_locked
			dll_delayctrl             : out   std_logic_vector(5 downto 0)                       -- dll_delayctrl
		);
	end component MebX_Qsys_Project_m2_ddr2_memory;

	component MebX_Qsys_Project_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(31 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component MebX_Qsys_Project_nios2_gen2_0;

	component MebX_Qsys_Project_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component MebX_Qsys_Project_onchip_memory;

	component MebX_Qsys_Project_pio_BUTTON is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component MebX_Qsys_Project_pio_BUTTON;

	component MebX_Qsys_Project_pio_DIP is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component MebX_Qsys_Project_pio_DIP;

	component MebX_Qsys_Project_pio_EXT is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_pio_EXT;

	component MebX_Qsys_Project_pio_LED is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_pio_LED;

	component MebX_Qsys_Project_pio_LED_painel is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(20 downto 0)                     -- export
		);
	end component MebX_Qsys_Project_pio_LED_painel;

	component MebX_Qsys_Project_pio_ctrl_io_lvds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_pio_ctrl_io_lvds;

	component MebX_Qsys_Project_pio_spw_demux_ch_1_select is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_pio_spw_demux_ch_1_select;

	component farm_rmap_memory_ffee_aeb_area_top is
		port (
			reset_i                     : in  std_logic                     := 'X';             -- reset
			clk_100_i                   : in  std_logic                     := 'X';             -- clk
			avs_rmap_0_address_i        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			avs_rmap_0_write_i          : in  std_logic                     := 'X';             -- write
			avs_rmap_0_read_i           : in  std_logic                     := 'X';             -- read
			avs_rmap_0_readdata_o       : out std_logic_vector(31 downto 0);                    -- readdata
			avs_rmap_0_writedata_i      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_rmap_0_waitrequest_o    : out std_logic;                                        -- waitrequest
			rms_rmap_0_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_0_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_0_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_0_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_0_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_0_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_0_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_0_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_1_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_1_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_1_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_1_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_1_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_1_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_1_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_1_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_2_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_2_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_2_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_2_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_2_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_2_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_2_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_2_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_3_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_3_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_3_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_3_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_3_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_3_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_3_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_3_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_4_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_4_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_4_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_4_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_4_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_4_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_4_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_4_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_5_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_5_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_5_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_5_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_5_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_5_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_5_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_5_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_6_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_6_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_6_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_6_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_6_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_6_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_6_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_6_rd_waitrequest_o : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_7_wr_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_7_write_i          : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_7_writedata_i      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_7_rd_address_i     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_7_read_i           : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_7_wr_waitrequest_o : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_7_readdata_o       : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_7_rd_waitrequest_o : out std_logic                                         -- rd_waitrequest_signal
		);
	end component farm_rmap_memory_ffee_aeb_area_top;

	component fdrm_rmap_memory_ffee_deb_area_top is
		port (
			reset_i                                  : in  std_logic                     := 'X';             -- reset
			clk_100_i                                : in  std_logic                     := 'X';             -- clk
			avs_rmap_0_address_i                     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			avs_rmap_0_write_i                       : in  std_logic                     := 'X';             -- write
			avs_rmap_0_read_i                        : in  std_logic                     := 'X';             -- read
			avs_rmap_0_readdata_o                    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_rmap_0_writedata_i                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_rmap_0_waitrequest_o                 : out std_logic;                                        -- waitrequest
			rms_rmap_0_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_0_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_0_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_0_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_0_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_0_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_0_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_0_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_1_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_1_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_1_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_1_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_1_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_1_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_1_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_1_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_2_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_2_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_2_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_2_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_2_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_2_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_2_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_2_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_3_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_3_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_3_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_3_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_3_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_3_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_3_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_3_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_4_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_4_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_4_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_4_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_4_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_4_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_4_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_4_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_5_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_5_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_5_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_5_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_5_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_5_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_5_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_5_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_6_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_6_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_6_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_6_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_6_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_6_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_6_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_6_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			rms_rmap_7_wr_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			rms_rmap_7_write_i                       : in  std_logic                     := 'X';             -- write_signal
			rms_rmap_7_writedata_i                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			rms_rmap_7_rd_address_i                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			rms_rmap_7_read_i                        : in  std_logic                     := 'X';             -- read_signal
			rms_rmap_7_wr_waitrequest_o              : out std_logic;                                        -- wr_waitrequest_signal
			rms_rmap_7_readdata_o                    : out std_logic_vector(7 downto 0);                     -- readdata_signal
			rms_rmap_7_rd_waitrequest_o              : out std_logic;                                        -- rd_waitrequest_signal
			avm_rmap_readdata_i                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			avm_rmap_waitrequest_i                   : in  std_logic                     := 'X';             -- waitrequest
			avm_rmap_address_o                       : out std_logic_vector(63 downto 0);                    -- address
			avm_rmap_read_o                          : out std_logic;                                        -- read
			avm_rmap_write_o                         : out std_logic;                                        -- write
			avm_rmap_writedata_o                     : out std_logic_vector(7 downto 0);                     -- writedata
			channel_hk_0_rmap_target_status_i        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rmap_target_status_signal
			channel_hk_0_rmap_target_indicate_i      : in  std_logic                     := 'X';             -- rmap_target_indicate_signal
			channel_hk_0_spw_link_escape_err_i       : in  std_logic                     := 'X';             -- spw_link_escape_err_signal
			channel_hk_0_spw_link_credit_err_i       : in  std_logic                     := 'X';             -- spw_link_credit_err_signal
			channel_hk_0_spw_link_parity_err_i       : in  std_logic                     := 'X';             -- spw_link_parity_err_signal
			channel_hk_0_spw_link_disconnect_i       : in  std_logic                     := 'X';             -- spw_link_disconnect_signal
			channel_hk_0_spw_link_started_i          : in  std_logic                     := 'X';             -- spw_link_started_signal
			channel_hk_0_spw_link_connecting_i       : in  std_logic                     := 'X';             -- spw_link_connecting_signal
			channel_hk_0_spw_link_running_i          : in  std_logic                     := 'X';             -- spw_link_running_signal
			channel_hk_0_frame_counter_i             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- frame_counter_signal
			channel_hk_0_left_buffer_ccd_number_i    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- left_buffer_ccd_number_signal
			channel_hk_0_right_buffer_ccd_number_i   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- right_buffer_ccd_number_signal
			channel_hk_0_left_buffer_ccd_side_i      : in  std_logic                     := 'X';             -- left_buffer_ccd_side_signal
			channel_hk_0_right_buffer_ccd_side_i     : in  std_logic                     := 'X';             -- right_buffer_ccd_side_signal
			channel_hk_0_err_left_buffer_overflow_i  : in  std_logic                     := 'X';             -- err_left_buffer_overflow_signal
			channel_hk_0_err_right_buffer_overflow_i : in  std_logic                     := 'X';             -- err_right_buffer_overflow_signal
			channel_hk_1_rmap_target_status_i        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rmap_target_status_signal
			channel_hk_1_rmap_target_indicate_i      : in  std_logic                     := 'X';             -- rmap_target_indicate_signal
			channel_hk_1_spw_link_escape_err_i       : in  std_logic                     := 'X';             -- spw_link_escape_err_signal
			channel_hk_1_spw_link_credit_err_i       : in  std_logic                     := 'X';             -- spw_link_credit_err_signal
			channel_hk_1_spw_link_parity_err_i       : in  std_logic                     := 'X';             -- spw_link_parity_err_signal
			channel_hk_1_spw_link_disconnect_i       : in  std_logic                     := 'X';             -- spw_link_disconnect_signal
			channel_hk_1_spw_link_started_i          : in  std_logic                     := 'X';             -- spw_link_started_signal
			channel_hk_1_spw_link_connecting_i       : in  std_logic                     := 'X';             -- spw_link_connecting_signal
			channel_hk_1_spw_link_running_i          : in  std_logic                     := 'X';             -- spw_link_running_signal
			channel_hk_1_frame_counter_i             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- frame_counter_signal
			channel_hk_1_left_buffer_ccd_number_i    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- left_buffer_ccd_number_signal
			channel_hk_1_right_buffer_ccd_number_i   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- right_buffer_ccd_number_signal
			channel_hk_1_left_buffer_ccd_side_i      : in  std_logic                     := 'X';             -- left_buffer_ccd_side_signal
			channel_hk_1_right_buffer_ccd_side_i     : in  std_logic                     := 'X';             -- right_buffer_ccd_side_signal
			channel_hk_1_err_left_buffer_overflow_i  : in  std_logic                     := 'X';             -- err_left_buffer_overflow_signal
			channel_hk_1_err_right_buffer_overflow_i : in  std_logic                     := 'X';             -- err_right_buffer_overflow_signal
			channel_hk_2_rmap_target_status_i        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rmap_target_status_signal
			channel_hk_2_rmap_target_indicate_i      : in  std_logic                     := 'X';             -- rmap_target_indicate_signal
			channel_hk_2_spw_link_escape_err_i       : in  std_logic                     := 'X';             -- spw_link_escape_err_signal
			channel_hk_2_spw_link_credit_err_i       : in  std_logic                     := 'X';             -- spw_link_credit_err_signal
			channel_hk_2_spw_link_parity_err_i       : in  std_logic                     := 'X';             -- spw_link_parity_err_signal
			channel_hk_2_spw_link_disconnect_i       : in  std_logic                     := 'X';             -- spw_link_disconnect_signal
			channel_hk_2_spw_link_started_i          : in  std_logic                     := 'X';             -- spw_link_started_signal
			channel_hk_2_spw_link_connecting_i       : in  std_logic                     := 'X';             -- spw_link_connecting_signal
			channel_hk_2_spw_link_running_i          : in  std_logic                     := 'X';             -- spw_link_running_signal
			channel_hk_2_frame_counter_i             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- frame_counter_signal
			channel_hk_2_left_buffer_ccd_number_i    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- left_buffer_ccd_number_signal
			channel_hk_2_right_buffer_ccd_number_i   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- right_buffer_ccd_number_signal
			channel_hk_2_left_buffer_ccd_side_i      : in  std_logic                     := 'X';             -- left_buffer_ccd_side_signal
			channel_hk_2_right_buffer_ccd_side_i     : in  std_logic                     := 'X';             -- right_buffer_ccd_side_signal
			channel_hk_2_err_left_buffer_overflow_i  : in  std_logic                     := 'X';             -- err_left_buffer_overflow_signal
			channel_hk_2_err_right_buffer_overflow_i : in  std_logic                     := 'X';             -- err_right_buffer_overflow_signal
			channel_hk_3_rmap_target_status_i        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rmap_target_status_signal
			channel_hk_3_rmap_target_indicate_i      : in  std_logic                     := 'X';             -- rmap_target_indicate_signal
			channel_hk_3_spw_link_escape_err_i       : in  std_logic                     := 'X';             -- spw_link_escape_err_signal
			channel_hk_3_spw_link_credit_err_i       : in  std_logic                     := 'X';             -- spw_link_credit_err_signal
			channel_hk_3_spw_link_parity_err_i       : in  std_logic                     := 'X';             -- spw_link_parity_err_signal
			channel_hk_3_spw_link_disconnect_i       : in  std_logic                     := 'X';             -- spw_link_disconnect_signal
			channel_hk_3_spw_link_started_i          : in  std_logic                     := 'X';             -- spw_link_started_signal
			channel_hk_3_spw_link_connecting_i       : in  std_logic                     := 'X';             -- spw_link_connecting_signal
			channel_hk_3_spw_link_running_i          : in  std_logic                     := 'X';             -- spw_link_running_signal
			channel_hk_3_frame_counter_i             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- frame_counter_signal
			channel_hk_3_left_buffer_ccd_number_i    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- left_buffer_ccd_number_signal
			channel_hk_3_right_buffer_ccd_number_i   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- right_buffer_ccd_number_signal
			channel_hk_3_left_buffer_ccd_side_i      : in  std_logic                     := 'X';             -- left_buffer_ccd_side_signal
			channel_hk_3_right_buffer_ccd_side_i     : in  std_logic                     := 'X';             -- right_buffer_ccd_side_signal
			channel_hk_3_err_left_buffer_overflow_i  : in  std_logic                     := 'X';             -- err_left_buffer_overflow_signal
			channel_hk_3_err_right_buffer_overflow_i : in  std_logic                     := 'X';             -- err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_i            : in  std_logic_vector(63 downto 0) := (others => 'X')  -- win_mem_addr_offset_signal
		);
	end component fdrm_rmap_memory_ffee_deb_area_top;

	component MebX_Qsys_Project_rs232_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_rs232_uart;

	component rst_controller_top is
		port (
			clock_sink_clk                          : in  std_logic                     := 'X';             -- clk
			reset_sink_reset                        : in  std_logic                     := 'X';             -- reset
			reset_source_rs232_reset                : out std_logic;                                        -- reset
			avalon_slave_rst_controller_address     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avalon_slave_rst_controller_write       : in  std_logic                     := 'X';             -- write
			avalon_slave_rst_controller_read        : in  std_logic                     := 'X';             -- read
			avalon_slave_rst_controller_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_rst_controller_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_rst_controller_waitrequest : out std_logic;                                        -- waitrequest
			simucam_reset_signal                    : out std_logic;                                        -- t_simucam_reset_signal
			reset_input_signal                      : in  std_logic                     := 'X'              -- t_reset_input_signal
		);
	end component rst_controller_top;

	component sync_ent is
		generic (
			g_SYNC_IRQ_NUMBER     : natural := 0;
			g_PRE_SYNC_IRQ_NUMBER : natural := 0
		);
		port (
			clock_sink_clk_i                 : in  std_logic                     := 'X';             -- clk
			reset_sink_reset_i               : in  std_logic                     := 'X';             -- reset
			avalon_slave_address_i           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avalon_slave_read_i              : in  std_logic                     := 'X';             -- read
			avalon_slave_write_i             : in  std_logic                     := 'X';             -- write
			avalon_slave_writedata_i         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_readdata_o          : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_waitrequest_o       : out std_logic;                                        -- waitrequest
			conduit_sync_signal_syncin_en_i  : in  std_logic                     := 'X';             -- conduit
			conduit_sync_signal_syncout_en_i : in  std_logic                     := 'X';             -- conduit
			conduit_sync_signal_syncin_i     : in  std_logic                     := 'X';             -- conduit
			conduit_sync_signal_spw1_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw2_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw3_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw4_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw5_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw6_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw7_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_spw8_o       : out std_logic;                                        -- conduit
			conduit_sync_signal_syncout_o    : out std_logic;                                        -- conduit
			sync_interrupt_sender_irq_o      : out std_logic;                                        -- irq
			pre_sync_interrupt_sender_irq_o  : out std_logic                                         -- irq
		);
	end component sync_ent;

	component MebX_Qsys_Project_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component MebX_Qsys_Project_sysid_qsys;

	component MebX_Qsys_Project_timer_1ms is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1ms;

	component MebX_Qsys_Project_timer_1us is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1us;

	component MebX_Qsys_Project_tristate_conduit_bridge_0 is
		port (
			clk                      : in    std_logic                     := 'X';             -- clk
			reset                    : in    std_logic                     := 'X';             -- reset
			request                  : in    std_logic                     := 'X';             -- request
			grant                    : out   std_logic;                                        -- grant
			tcs_tcm_address_out      : in    std_logic_vector(25 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out         : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen       : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in          : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out          : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tcm_read_n_out           : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component MebX_Qsys_Project_tristate_conduit_bridge_0;

	component MebX_Qsys_Project_mm_interconnect_0 is
		port (
			clk_100_clk_clk                                                       : in  std_logic                      := 'X';             -- clk
			m2_ddr2_memory_afi_clk_clk                                            : in  std_logic                      := 'X';             -- clk
			m2_ddr2_memory_afi_half_clk_clk                                       : in  std_logic                      := 'X';             -- clk
			FTDI_UMFT601A_Module_reset_sink_reset_bridge_in_reset_reset           : in  std_logic                      := 'X';             -- reset
			m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset                  : in  std_logic                      := 'X';             -- reset
			m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset       : in  std_logic                      := 'X';             -- reset
			m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset                 : in  std_logic                      := 'X';             -- reset
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_address      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_waitrequest  : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_read         : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_readdata     : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_address     : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_waitrequest : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_read        : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_readdata    : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_address      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_waitrequest  : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_read         : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_readdata     : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_address     : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_waitrequest : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_read        : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_readdata    : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_address      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_waitrequest  : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_read         : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_readdata     : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_address     : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_waitrequest : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_read        : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_readdata    : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_address      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_waitrequest  : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_read         : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_readdata     : out std_logic_vector(255 downto 0);                    -- readdata
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_address     : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_waitrequest : out std_logic;                                         -- waitrequest
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_read        : in  std_logic                      := 'X';             -- read
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_readdata    : out std_logic_vector(255 downto 0);                    -- readdata
			ddr2_address_span_extender_expanded_master_address                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			ddr2_address_span_extender_expanded_master_waitrequest                : out std_logic;                                         -- waitrequest
			ddr2_address_span_extender_expanded_master_burstcount                 : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			ddr2_address_span_extender_expanded_master_byteenable                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			ddr2_address_span_extender_expanded_master_read                       : in  std_logic                      := 'X';             -- read
			ddr2_address_span_extender_expanded_master_readdata                   : out std_logic_vector(31 downto 0);                     -- readdata
			ddr2_address_span_extender_expanded_master_readdatavalid              : out std_logic;                                         -- readdatavalid
			ddr2_address_span_extender_expanded_master_write                      : in  std_logic                      := 'X';             -- write
			ddr2_address_span_extender_expanded_master_writedata                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			FTDI_UMFT601A_Module_avalon_imgt_master_data_address                  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			FTDI_UMFT601A_Module_avalon_imgt_master_data_waitrequest              : out std_logic;                                         -- waitrequest
			FTDI_UMFT601A_Module_avalon_imgt_master_data_write                    : in  std_logic                      := 'X';             -- write
			FTDI_UMFT601A_Module_avalon_imgt_master_data_writedata                : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- writedata
			FTDI_UMFT601A_Module_avalon_master_data_address                       : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			FTDI_UMFT601A_Module_avalon_master_data_waitrequest                   : out std_logic;                                         -- waitrequest
			FTDI_UMFT601A_Module_avalon_master_data_read                          : in  std_logic                      := 'X';             -- read
			FTDI_UMFT601A_Module_avalon_master_data_readdata                      : out std_logic_vector(255 downto 0);                    -- readdata
			FTDI_UMFT601A_Module_avalon_master_data_write                         : in  std_logic                      := 'X';             -- write
			FTDI_UMFT601A_Module_avalon_master_data_writedata                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			Memory_Filler_avalon_master_data_address                              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Memory_Filler_avalon_master_data_waitrequest                          : out std_logic;                                         -- waitrequest
			Memory_Filler_avalon_master_data_write                                : in  std_logic                      := 'X';             -- write
			Memory_Filler_avalon_master_data_writedata                            : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address                  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest              : out std_logic;                                         -- waitrequest
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read                     : in  std_logic                      := 'X';             -- read
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata                 : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write                    : in  std_logic                      := 'X';             -- write
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			m1_clock_bridge_s0_address                                            : out std_logic_vector(30 downto 0);                     -- address
			m1_clock_bridge_s0_write                                              : out std_logic;                                         -- write
			m1_clock_bridge_s0_read                                               : out std_logic;                                         -- read
			m1_clock_bridge_s0_readdata                                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m1_clock_bridge_s0_writedata                                          : out std_logic_vector(255 downto 0);                    -- writedata
			m1_clock_bridge_s0_burstcount                                         : out std_logic_vector(2 downto 0);                      -- burstcount
			m1_clock_bridge_s0_byteenable                                         : out std_logic_vector(31 downto 0);                     -- byteenable
			m1_clock_bridge_s0_readdatavalid                                      : in  std_logic                      := 'X';             -- readdatavalid
			m1_clock_bridge_s0_waitrequest                                        : in  std_logic                      := 'X';             -- waitrequest
			m1_clock_bridge_s0_debugaccess                                        : out std_logic;                                         -- debugaccess
			m2_ddr2_memory_avl_address                                            : out std_logic_vector(25 downto 0);                     -- address
			m2_ddr2_memory_avl_write                                              : out std_logic;                                         -- write
			m2_ddr2_memory_avl_read                                               : out std_logic;                                         -- read
			m2_ddr2_memory_avl_readdata                                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_memory_avl_writedata                                          : out std_logic_vector(255 downto 0);                    -- writedata
			m2_ddr2_memory_avl_beginbursttransfer                                 : out std_logic;                                         -- beginbursttransfer
			m2_ddr2_memory_avl_burstcount                                         : out std_logic_vector(7 downto 0);                      -- burstcount
			m2_ddr2_memory_avl_byteenable                                         : out std_logic_vector(31 downto 0);                     -- byteenable
			m2_ddr2_memory_avl_readdatavalid                                      : in  std_logic                      := 'X';             -- readdatavalid
			m2_ddr2_memory_avl_waitrequest                                        : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_0;

	component MebX_Qsys_Project_mm_interconnect_1 is
		port (
			clk_100_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			ext_flash_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_burstcount                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			nios2_gen2_0_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			clock_bridge_afi_50_s0_address                                 : out std_logic_vector(11 downto 0);                    -- address
			clock_bridge_afi_50_s0_write                                   : out std_logic;                                        -- write
			clock_bridge_afi_50_s0_read                                    : out std_logic;                                        -- read
			clock_bridge_afi_50_s0_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clock_bridge_afi_50_s0_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			clock_bridge_afi_50_s0_burstcount                              : out std_logic_vector(0 downto 0);                     -- burstcount
			clock_bridge_afi_50_s0_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			clock_bridge_afi_50_s0_readdatavalid                           : in  std_logic                     := 'X';             -- readdatavalid
			clock_bridge_afi_50_s0_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			clock_bridge_afi_50_s0_debugaccess                             : out std_logic;                                        -- debugaccess
			Communication_Module_v2_Ch1_avalon_mm_config_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Communication_Module_v2_Ch1_avalon_mm_config_slave_write       : out std_logic;                                        -- write
			Communication_Module_v2_Ch1_avalon_mm_config_slave_read        : out std_logic;                                        -- read
			Communication_Module_v2_Ch1_avalon_mm_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Communication_Module_v2_Ch1_avalon_mm_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Communication_Module_v2_Ch1_avalon_mm_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			Communication_Module_v2_Ch2_avalon_mm_config_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Communication_Module_v2_Ch2_avalon_mm_config_slave_write       : out std_logic;                                        -- write
			Communication_Module_v2_Ch2_avalon_mm_config_slave_read        : out std_logic;                                        -- read
			Communication_Module_v2_Ch2_avalon_mm_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Communication_Module_v2_Ch2_avalon_mm_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Communication_Module_v2_Ch2_avalon_mm_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			Communication_Module_v2_Ch3_avalon_mm_config_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Communication_Module_v2_Ch3_avalon_mm_config_slave_write       : out std_logic;                                        -- write
			Communication_Module_v2_Ch3_avalon_mm_config_slave_read        : out std_logic;                                        -- read
			Communication_Module_v2_Ch3_avalon_mm_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Communication_Module_v2_Ch3_avalon_mm_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Communication_Module_v2_Ch3_avalon_mm_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			Communication_Module_v2_Ch4_avalon_mm_config_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Communication_Module_v2_Ch4_avalon_mm_config_slave_write       : out std_logic;                                        -- write
			Communication_Module_v2_Ch4_avalon_mm_config_slave_read        : out std_logic;                                        -- read
			Communication_Module_v2_Ch4_avalon_mm_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Communication_Module_v2_Ch4_avalon_mm_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Communication_Module_v2_Ch4_avalon_mm_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			ddr2_address_span_extender_cntl_write                          : out std_logic;                                        -- write
			ddr2_address_span_extender_cntl_read                           : out std_logic;                                        -- read
			ddr2_address_span_extender_cntl_readdata                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			ddr2_address_span_extender_cntl_writedata                      : out std_logic_vector(63 downto 0);                    -- writedata
			ddr2_address_span_extender_cntl_byteenable                     : out std_logic_vector(7 downto 0);                     -- byteenable
			ddr2_address_span_extender_windowed_slave_address              : out std_logic_vector(28 downto 0);                    -- address
			ddr2_address_span_extender_windowed_slave_write                : out std_logic;                                        -- write
			ddr2_address_span_extender_windowed_slave_read                 : out std_logic;                                        -- read
			ddr2_address_span_extender_windowed_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ddr2_address_span_extender_windowed_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			ddr2_address_span_extender_windowed_slave_burstcount           : out std_logic_vector(7 downto 0);                     -- burstcount
			ddr2_address_span_extender_windowed_slave_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			ext_flash_uas_address                                          : out std_logic_vector(25 downto 0);                    -- address
			ext_flash_uas_write                                            : out std_logic;                                        -- write
			ext_flash_uas_read                                             : out std_logic;                                        -- read
			ext_flash_uas_readdata                                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			ext_flash_uas_writedata                                        : out std_logic_vector(15 downto 0);                    -- writedata
			ext_flash_uas_burstcount                                       : out std_logic_vector(1 downto 0);                     -- burstcount
			ext_flash_uas_byteenable                                       : out std_logic_vector(1 downto 0);                     -- byteenable
			ext_flash_uas_readdatavalid                                    : in  std_logic                     := 'X';             -- readdatavalid
			ext_flash_uas_waitrequest                                      : in  std_logic                     := 'X';             -- waitrequest
			ext_flash_uas_lock                                             : out std_logic;                                        -- lock
			ext_flash_uas_debugaccess                                      : out std_logic;                                        -- debugaccess
			FTDI_UMFT601A_Module_avalon_slave_config_address               : out std_logic_vector(7 downto 0);                     -- address
			FTDI_UMFT601A_Module_avalon_slave_config_write                 : out std_logic;                                        -- write
			FTDI_UMFT601A_Module_avalon_slave_config_read                  : out std_logic;                                        -- read
			FTDI_UMFT601A_Module_avalon_slave_config_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			FTDI_UMFT601A_Module_avalon_slave_config_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			FTDI_UMFT601A_Module_avalon_slave_config_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                       : out std_logic;                                        -- chipselect
			Memory_Filler_avalon_slave_config_address                      : out std_logic_vector(7 downto 0);                     -- address
			Memory_Filler_avalon_slave_config_write                        : out std_logic;                                        -- write
			Memory_Filler_avalon_slave_config_read                         : out std_logic;                                        -- read
			Memory_Filler_avalon_slave_config_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Memory_Filler_avalon_slave_config_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			Memory_Filler_avalon_slave_config_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Memory_Filler_avalon_slave_config_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                                       : out std_logic_vector(17 downto 0);                    -- address
			onchip_memory_s1_write                                         : out std_logic;                                        -- write
			onchip_memory_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                                    : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                                    : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                                         : out std_logic;                                        -- clken
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address           : out std_logic_vector(11 downto 0);                    -- address
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write             : out std_logic;                                        -- write
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read              : out std_logic;                                        -- read
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address           : out std_logic_vector(11 downto 0);                    -- address
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write             : out std_logic;                                        -- write
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read              : out std_logic;                                        -- read
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address           : out std_logic_vector(11 downto 0);                    -- address
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write             : out std_logic;                                        -- write
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read              : out std_logic;                                        -- read
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address           : out std_logic_vector(11 downto 0);                    -- address
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write             : out std_logic;                                        -- write
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read              : out std_logic;                                        -- read
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address             : out std_logic_vector(11 downto 0);                    -- address
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write               : out std_logic;                                        -- write
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read                : out std_logic;                                        -- read
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			sysid_qsys_control_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component MebX_Qsys_Project_mm_interconnect_1;

	component MebX_Qsys_Project_mm_interconnect_2 is
		port (
			clk_50_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			rs232_uart_reset_reset_bridge_in_reset_reset                         : in  std_logic                     := 'X';             -- reset
			clock_bridge_afi_50_m0_address                                       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_bridge_afi_50_m0_waitrequest                                   : out std_logic;                                        -- waitrequest
			clock_bridge_afi_50_m0_burstcount                                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_bridge_afi_50_m0_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_bridge_afi_50_m0_read                                          : in  std_logic                     := 'X';             -- read
			clock_bridge_afi_50_m0_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			clock_bridge_afi_50_m0_readdatavalid                                 : out std_logic;                                        -- readdatavalid
			clock_bridge_afi_50_m0_write                                         : in  std_logic                     := 'X';             -- write
			clock_bridge_afi_50_m0_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_bridge_afi_50_m0_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     : out std_logic_vector(7 downto 0);                     -- address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       : out std_logic;                                        -- write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        : out std_logic;                                        -- read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  : out std_logic;                                        -- chipselect
			csense_adc_fo_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			csense_adc_fo_s1_write                                               : out std_logic;                                        -- write
			csense_adc_fo_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_adc_fo_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			csense_adc_fo_s1_chipselect                                          : out std_logic;                                        -- chipselect
			csense_cs_n_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			csense_cs_n_s1_write                                                 : out std_logic;                                        -- write
			csense_cs_n_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_cs_n_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			csense_cs_n_s1_chipselect                                            : out std_logic;                                        -- chipselect
			csense_sck_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			csense_sck_s1_write                                                  : out std_logic;                                        -- write
			csense_sck_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sck_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sck_s1_chipselect                                             : out std_logic;                                        -- chipselect
			csense_sdi_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			csense_sdi_s1_write                                                  : out std_logic;                                        -- write
			csense_sdi_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sdi_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sdi_s1_chipselect                                             : out std_logic;                                        -- chipselect
			csense_sdo_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			csense_sdo_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_scl_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			m1_ddr2_i2c_scl_s1_write                                             : out std_logic;                                        -- write
			m1_ddr2_i2c_scl_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_scl_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			m1_ddr2_i2c_scl_s1_chipselect                                        : out std_logic;                                        -- chipselect
			m1_ddr2_i2c_sda_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			m1_ddr2_i2c_sda_s1_write                                             : out std_logic;                                        -- write
			m1_ddr2_i2c_sda_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_sda_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			m1_ddr2_i2c_sda_s1_chipselect                                        : out std_logic;                                        -- chipselect
			m2_ddr2_i2c_scl_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			m2_ddr2_i2c_scl_s1_write                                             : out std_logic;                                        -- write
			m2_ddr2_i2c_scl_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_i2c_scl_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			m2_ddr2_i2c_scl_s1_chipselect                                        : out std_logic;                                        -- chipselect
			m2_ddr2_i2c_sda_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			m2_ddr2_i2c_sda_s1_write                                             : out std_logic;                                        -- write
			m2_ddr2_i2c_sda_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_i2c_sda_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			m2_ddr2_i2c_sda_s1_chipselect                                        : out std_logic;                                        -- chipselect
			pio_BUTTON_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			pio_BUTTON_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ctrl_io_lvds_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			pio_ctrl_io_lvds_s1_write                                            : out std_logic;                                        -- write
			pio_ctrl_io_lvds_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ctrl_io_lvds_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			pio_ctrl_io_lvds_s1_chipselect                                       : out std_logic;                                        -- chipselect
			pio_DIP_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			pio_DIP_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_EXT_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			pio_EXT_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ftdi_umft601a_module_reset_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			pio_ftdi_umft601a_module_reset_s1_write                              : out std_logic;                                        -- write
			pio_ftdi_umft601a_module_reset_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ftdi_umft601a_module_reset_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_ftdi_umft601a_module_reset_s1_chipselect                         : out std_logic;                                        -- chipselect
			pio_iso_logic_signal_enable_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pio_iso_logic_signal_enable_s1_write                                 : out std_logic;                                        -- write
			pio_iso_logic_signal_enable_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_iso_logic_signal_enable_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_iso_logic_signal_enable_s1_chipselect                            : out std_logic;                                        -- chipselect
			pio_LED_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			pio_LED_s1_write                                                     : out std_logic;                                        -- write
			pio_LED_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_LED_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			pio_LED_s1_chipselect                                                : out std_logic;                                        -- chipselect
			pio_LED_painel_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			pio_LED_painel_s1_write                                              : out std_logic;                                        -- write
			pio_LED_painel_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_LED_painel_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_LED_painel_s1_chipselect                                         : out std_logic;                                        -- chipselect
			pio_spw_demux_ch_1_select_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_spw_demux_ch_1_select_s1_write                                   : out std_logic;                                        -- write
			pio_spw_demux_ch_1_select_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_spw_demux_ch_1_select_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_spw_demux_ch_1_select_s1_chipselect                              : out std_logic;                                        -- chipselect
			pio_spw_demux_ch_2_select_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_spw_demux_ch_2_select_s1_write                                   : out std_logic;                                        -- write
			pio_spw_demux_ch_2_select_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_spw_demux_ch_2_select_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_spw_demux_ch_2_select_s1_chipselect                              : out std_logic;                                        -- chipselect
			pio_spw_demux_ch_3_select_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_spw_demux_ch_3_select_s1_write                                   : out std_logic;                                        -- write
			pio_spw_demux_ch_3_select_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_spw_demux_ch_3_select_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_spw_demux_ch_3_select_s1_chipselect                              : out std_logic;                                        -- chipselect
			pio_spw_demux_ch_4_select_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_spw_demux_ch_4_select_s1_write                                   : out std_logic;                                        -- write
			pio_spw_demux_ch_4_select_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_spw_demux_ch_4_select_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_spw_demux_ch_4_select_s1_chipselect                              : out std_logic;                                        -- chipselect
			rs232_uart_s1_address                                                : out std_logic_vector(2 downto 0);                     -- address
			rs232_uart_s1_write                                                  : out std_logic;                                        -- write
			rs232_uart_s1_read                                                   : out std_logic;                                        -- read
			rs232_uart_s1_readdata                                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			rs232_uart_s1_writedata                                              : out std_logic_vector(15 downto 0);                    -- writedata
			rs232_uart_s1_begintransfer                                          : out std_logic;                                        -- begintransfer
			rs232_uart_s1_chipselect                                             : out std_logic;                                        -- chipselect
			rst_controller_avalon_rst_controller_slave_address                   : out std_logic_vector(3 downto 0);                     -- address
			rst_controller_avalon_rst_controller_slave_write                     : out std_logic;                                        -- write
			rst_controller_avalon_rst_controller_slave_read                      : out std_logic;                                        -- read
			rst_controller_avalon_rst_controller_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rst_controller_avalon_rst_controller_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			rst_controller_avalon_rst_controller_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			rtcc_alarm_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			rtcc_alarm_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_cs_n_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			rtcc_cs_n_s1_write                                                   : out std_logic;                                        -- write
			rtcc_cs_n_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_cs_n_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_cs_n_s1_chipselect                                              : out std_logic;                                        -- chipselect
			rtcc_sck_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sck_s1_write                                                    : out std_logic;                                        -- write
			rtcc_sck_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_sck_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_sck_s1_chipselect                                               : out std_logic;                                        -- chipselect
			rtcc_sdi_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sdi_s1_write                                                    : out std_logic;                                        -- write
			rtcc_sdi_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_sdi_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_sdi_s1_chipselect                                               : out std_logic;                                        -- chipselect
			rtcc_sdo_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sdo_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sd_card_wp_n_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			sd_card_wp_n_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sync_avalon_mm_slave_address                                         : out std_logic_vector(7 downto 0);                     -- address
			sync_avalon_mm_slave_write                                           : out std_logic;                                        -- write
			sync_avalon_mm_slave_read                                            : out std_logic;                                        -- read
			sync_avalon_mm_slave_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sync_avalon_mm_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			sync_avalon_mm_slave_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			temp_scl_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			temp_scl_s1_write                                                    : out std_logic;                                        -- write
			temp_scl_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_scl_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			temp_scl_s1_chipselect                                               : out std_logic;                                        -- chipselect
			temp_sda_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			temp_sda_s1_write                                                    : out std_logic;                                        -- write
			temp_sda_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_sda_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			temp_sda_s1_chipselect                                               : out std_logic;                                        -- chipselect
			timer_1ms_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			timer_1ms_s1_write                                                   : out std_logic;                                        -- write
			timer_1ms_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1ms_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1ms_s1_chipselect                                              : out std_logic;                                        -- chipselect
			timer_1us_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			timer_1us_s1_write                                                   : out std_logic;                                        -- write
			timer_1us_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1us_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1us_s1_chipselect                                              : out std_logic                                         -- chipselect
		);
	end component MebX_Qsys_Project_mm_interconnect_2;

	component MebX_Qsys_Project_mm_interconnect_3 is
		port (
			m1_ddr2_memory_afi_clk_clk                                      : in  std_logic                      := 'X';             -- clk
			m1_ddr2_memory_afi_half_clk_clk                                 : in  std_logic                      := 'X';             -- clk
			m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset            : in  std_logic                      := 'X';             -- reset
			m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           : in  std_logic                      := 'X';             -- reset
			m1_clock_bridge_m0_address                                      : in  std_logic_vector(30 downto 0)  := (others => 'X'); -- address
			m1_clock_bridge_m0_waitrequest                                  : out std_logic;                                         -- waitrequest
			m1_clock_bridge_m0_burstcount                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			m1_clock_bridge_m0_byteenable                                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			m1_clock_bridge_m0_read                                         : in  std_logic                      := 'X';             -- read
			m1_clock_bridge_m0_readdata                                     : out std_logic_vector(255 downto 0);                    -- readdata
			m1_clock_bridge_m0_readdatavalid                                : out std_logic;                                         -- readdatavalid
			m1_clock_bridge_m0_write                                        : in  std_logic                      := 'X';             -- write
			m1_clock_bridge_m0_writedata                                    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			m1_clock_bridge_m0_debugaccess                                  : in  std_logic                      := 'X';             -- debugaccess
			m1_ddr2_memory_avl_address                                      : out std_logic_vector(25 downto 0);                     -- address
			m1_ddr2_memory_avl_write                                        : out std_logic;                                         -- write
			m1_ddr2_memory_avl_read                                         : out std_logic;                                         -- read
			m1_ddr2_memory_avl_readdata                                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_memory_avl_writedata                                    : out std_logic_vector(255 downto 0);                    -- writedata
			m1_ddr2_memory_avl_beginbursttransfer                           : out std_logic;                                         -- beginbursttransfer
			m1_ddr2_memory_avl_burstcount                                   : out std_logic_vector(7 downto 0);                      -- burstcount
			m1_ddr2_memory_avl_byteenable                                   : out std_logic_vector(31 downto 0);                     -- byteenable
			m1_ddr2_memory_avl_readdatavalid                                : in  std_logic                      := 'X';             -- readdatavalid
			m1_ddr2_memory_avl_waitrequest                                  : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_3;

	component MebX_Qsys_Project_irq_mapper is
		port (
			clk            : in  std_logic                     := 'X'; -- clk
			reset          : in  std_logic                     := 'X'; -- reset
			receiver0_irq  : in  std_logic                     := 'X'; -- irq
			receiver1_irq  : in  std_logic                     := 'X'; -- irq
			receiver2_irq  : in  std_logic                     := 'X'; -- irq
			receiver3_irq  : in  std_logic                     := 'X'; -- irq
			receiver4_irq  : in  std_logic                     := 'X'; -- irq
			receiver5_irq  : in  std_logic                     := 'X'; -- irq
			receiver6_irq  : in  std_logic                     := 'X'; -- irq
			receiver7_irq  : in  std_logic                     := 'X'; -- irq
			receiver8_irq  : in  std_logic                     := 'X'; -- irq
			receiver9_irq  : in  std_logic                     := 'X'; -- irq
			receiver10_irq : in  std_logic                     := 'X'; -- irq
			receiver11_irq : in  std_logic                     := 'X'; -- irq
			receiver12_irq : in  std_logic                     := 'X'; -- irq
			receiver13_irq : in  std_logic                     := 'X'; -- irq
			receiver14_irq : in  std_logic                     := 'X'; -- irq
			receiver15_irq : in  std_logic                     := 'X'; -- irq
			sender_irq     : out std_logic_vector(31 downto 0)         -- irq
		);
	end component MebX_Qsys_Project_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component mebx_qsys_project_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_001;

	component mebx_qsys_project_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_002;

	component mebx_qsys_project_rst_controller_004 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_004;

	component mebx_qsys_project_clock_bridge_afi_50 is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             --   m0_clk.clk
			m0_reset         : in  std_logic                     := 'X';             -- m0_reset.reset
			s0_clk           : in  std_logic                     := 'X';             --   s0_clk.clk
			s0_reset         : in  std_logic                     := 'X';             -- s0_reset.reset
			s0_waitrequest   : out std_logic;                                        --       s0.waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    --         .readdata
			s0_readdatavalid : out std_logic;                                        --         .readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); --         .burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); --         .writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); --         .address
			s0_write         : in  std_logic                     := 'X';             --         .write
			s0_read          : in  std_logic                     := 'X';             --         .read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); --         .byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             --         .debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             --       m0.waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); --         .readdata
			m0_readdatavalid : in  std_logic                     := 'X';             --         .readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     --         .burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    --         .writedata
			m0_address       : out std_logic_vector(11 downto 0);                    --         .address
			m0_write         : out std_logic;                                        --         .write
			m0_read          : out std_logic;                                        --         .read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     --         .byteenable
			m0_debugaccess   : out std_logic                                         --         .debugaccess
		);
	end component mebx_qsys_project_clock_bridge_afi_50;

	component mebx_qsys_project_m1_clock_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                      := 'X';             --   m0_clk.clk
			m0_reset         : in  std_logic                      := 'X';             -- m0_reset.reset
			s0_clk           : in  std_logic                      := 'X';             --   s0_clk.clk
			s0_reset         : in  std_logic                      := 'X';             -- s0_reset.reset
			s0_waitrequest   : out std_logic;                                         --       s0.waitrequest
			s0_readdata      : out std_logic_vector(255 downto 0);                    --         .readdata
			s0_readdatavalid : out std_logic;                                         --         .readdatavalid
			s0_burstcount    : in  std_logic_vector(2 downto 0)   := (others => 'X'); --         .burstcount
			s0_writedata     : in  std_logic_vector(255 downto 0) := (others => 'X'); --         .writedata
			s0_address       : in  std_logic_vector(30 downto 0)  := (others => 'X'); --         .address
			s0_write         : in  std_logic                      := 'X';             --         .write
			s0_read          : in  std_logic                      := 'X';             --         .read
			s0_byteenable    : in  std_logic_vector(31 downto 0)  := (others => 'X'); --         .byteenable
			s0_debugaccess   : in  std_logic                      := 'X';             --         .debugaccess
			m0_waitrequest   : in  std_logic                      := 'X';             --       m0.waitrequest
			m0_readdata      : in  std_logic_vector(255 downto 0) := (others => 'X'); --         .readdata
			m0_readdatavalid : in  std_logic                      := 'X';             --         .readdatavalid
			m0_burstcount    : out std_logic_vector(2 downto 0);                      --         .burstcount
			m0_writedata     : out std_logic_vector(255 downto 0);                    --         .writedata
			m0_address       : out std_logic_vector(30 downto 0);                     --         .address
			m0_write         : out std_logic;                                         --         .write
			m0_read          : out std_logic;                                         --         .read
			m0_byteenable    : out std_logic_vector(31 downto 0);                     --         .byteenable
			m0_debugaccess   : out std_logic                                          --         .debugaccess
		);
	end component mebx_qsys_project_m1_clock_bridge;

	signal m2_ddr2_memory_afi_clk_clk                                                                       : std_logic;                      -- m2_ddr2_memory:afi_clk -> [SpaceWire_Channel_A:clk_200_i, SpaceWire_Channel_B:clk_200_i, SpaceWire_Channel_C:clk_200_i, SpaceWire_Channel_D:clk_200_i, SpaceWire_Channel_E:clk_200_i, SpaceWire_Channel_F:clk_200_i, SpaceWire_Channel_G:clk_200_i, SpaceWire_Channel_H:clk_200_i, mm_interconnect_0:m2_ddr2_memory_afi_clk_clk, rst_controller_003:clk]
	signal m2_ddr2_memory_afi_half_clk_clk                                                                  : std_logic;                      -- m2_ddr2_memory:afi_half_clk -> [Communication_Module_v2_Ch1:clock_sink_clk_i, Communication_Module_v2_Ch2:clock_sink_clk_i, Communication_Module_v2_Ch3:clock_sink_clk_i, Communication_Module_v2_Ch4:clock_sink_clk_i, FTDI_UMFT601A_Module:clock_sink_clk_i, Memory_Filler:clock_sink_clk_i, SpaceWire_Channel_A:clk_100_i, SpaceWire_Channel_B:clk_100_i, SpaceWire_Channel_C:clk_100_i, SpaceWire_Channel_D:clk_100_i, SpaceWire_Channel_E:clk_100_i, SpaceWire_Channel_F:clk_100_i, SpaceWire_Channel_G:clk_100_i, SpaceWire_Channel_H:clk_100_i, SpaceWire_Demux_Ch1:clock_i, SpaceWire_Demux_Ch2:clock_i, SpaceWire_Demux_Ch3:clock_i, SpaceWire_Demux_Ch4:clock_i, clock_bridge_afi_50:s0_clk, ddr2_address_span_extender:clk, ext_flash:clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, jtag_uart_0:clk, m1_clock_bridge:s0_clk, mm_interconnect_0:clk_100_clk_clk, mm_interconnect_0:m2_ddr2_memory_afi_half_clk_clk, mm_interconnect_1:clk_100_clk_clk, nios2_gen2_0:clk, onchip_memory:clk, rmap_mem_ffee_aeb_1_area:clk_100_i, rmap_mem_ffee_aeb_2_area:clk_100_i, rmap_mem_ffee_aeb_3_area:clk_100_i, rmap_mem_ffee_aeb_4_area:clk_100_i, rmap_mem_ffee_deb_area:clk_100_i, rst_controller_002:clk, rst_controller_004:clk, rst_controller_006:clk, sysid_qsys:clock, tristate_conduit_bridge_0:clk]
	signal m1_ddr2_memory_afi_half_clk_clk                                                                  : std_logic;                      -- m1_ddr2_memory:afi_half_clk -> [m1_clock_bridge:m0_clk, mm_interconnect_3:m1_ddr2_memory_afi_half_clk_clk, rst_controller_005:clk]
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_number_signal             : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch4:channel_hk_left_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_3_left_buffer_ccd_number_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_side_signal              : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_right_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_3_right_buffer_ccd_side_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_escape_err_signal                : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_escape_err_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_escape_err_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_indicate_signal               : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_rmap_target_indicate_o -> rmap_mem_ffee_deb_area:channel_hk_3_rmap_target_indicate_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_running_signal                   : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_running_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_running_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_credit_err_signal                : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_credit_err_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_credit_err_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_side_signal               : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_left_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_3_left_buffer_ccd_side_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_err_right_buffer_overflow_signal          : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_err_right_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_3_err_right_buffer_overflow_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_status_signal                 : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:channel_hk_rmap_target_status_o -> rmap_mem_ffee_deb_area:channel_hk_3_rmap_target_status_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_parity_err_signal                : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_parity_err_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_parity_err_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_disconnect_signal                : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_disconnect_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_disconnect_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_connecting_signal                : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_connecting_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_connecting_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_started_signal                   : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_spw_link_started_o -> rmap_mem_ffee_deb_area:channel_hk_3_spw_link_started_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_number_signal            : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch4:channel_hk_right_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_3_right_buffer_ccd_number_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_frame_counter_signal                      : std_logic_vector(15 downto 0);  -- Communication_Module_v2_Ch4:channel_hk_frame_counter_o -> rmap_mem_ffee_deb_area:channel_hk_3_frame_counter_i
	signal communication_module_v2_ch4_conduit_end_channel_hk_out_err_left_buffer_overflow_signal           : std_logic;                      -- Communication_Module_v2_Ch4:channel_hk_err_left_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_3_err_left_buffer_overflow_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_number_signal             : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch1:channel_hk_left_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_0_left_buffer_ccd_number_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_side_signal              : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_right_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_0_right_buffer_ccd_side_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_escape_err_signal                : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_escape_err_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_escape_err_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_indicate_signal               : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_rmap_target_indicate_o -> rmap_mem_ffee_deb_area:channel_hk_0_rmap_target_indicate_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_running_signal                   : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_running_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_running_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_credit_err_signal                : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_credit_err_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_credit_err_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_side_signal               : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_left_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_0_left_buffer_ccd_side_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_err_right_buffer_overflow_signal          : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_err_right_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_0_err_right_buffer_overflow_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_status_signal                 : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:channel_hk_rmap_target_status_o -> rmap_mem_ffee_deb_area:channel_hk_0_rmap_target_status_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_parity_err_signal                : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_parity_err_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_parity_err_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_disconnect_signal                : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_disconnect_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_disconnect_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_connecting_signal                : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_connecting_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_connecting_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_started_signal                   : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_spw_link_started_o -> rmap_mem_ffee_deb_area:channel_hk_0_spw_link_started_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_number_signal            : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch1:channel_hk_right_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_0_right_buffer_ccd_number_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_frame_counter_signal                      : std_logic_vector(15 downto 0);  -- Communication_Module_v2_Ch1:channel_hk_frame_counter_o -> rmap_mem_ffee_deb_area:channel_hk_0_frame_counter_i
	signal communication_module_v2_ch1_conduit_end_channel_hk_out_err_left_buffer_overflow_signal           : std_logic;                      -- Communication_Module_v2_Ch1:channel_hk_err_left_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_0_err_left_buffer_overflow_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_number_signal             : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch2:channel_hk_left_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_1_left_buffer_ccd_number_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_side_signal              : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_right_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_1_right_buffer_ccd_side_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_escape_err_signal                : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_escape_err_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_escape_err_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_indicate_signal               : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_rmap_target_indicate_o -> rmap_mem_ffee_deb_area:channel_hk_1_rmap_target_indicate_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_running_signal                   : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_running_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_running_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_credit_err_signal                : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_credit_err_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_credit_err_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_side_signal               : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_left_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_1_left_buffer_ccd_side_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_err_right_buffer_overflow_signal          : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_err_right_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_1_err_right_buffer_overflow_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_status_signal                 : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:channel_hk_rmap_target_status_o -> rmap_mem_ffee_deb_area:channel_hk_1_rmap_target_status_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_parity_err_signal                : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_parity_err_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_parity_err_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_disconnect_signal                : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_disconnect_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_disconnect_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_connecting_signal                : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_connecting_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_connecting_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_started_signal                   : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_spw_link_started_o -> rmap_mem_ffee_deb_area:channel_hk_1_spw_link_started_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_number_signal            : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch2:channel_hk_right_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_1_right_buffer_ccd_number_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_frame_counter_signal                      : std_logic_vector(15 downto 0);  -- Communication_Module_v2_Ch2:channel_hk_frame_counter_o -> rmap_mem_ffee_deb_area:channel_hk_1_frame_counter_i
	signal communication_module_v2_ch2_conduit_end_channel_hk_out_err_left_buffer_overflow_signal           : std_logic;                      -- Communication_Module_v2_Ch2:channel_hk_err_left_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_1_err_left_buffer_overflow_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_number_signal             : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch3:channel_hk_left_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_2_left_buffer_ccd_number_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_side_signal              : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_right_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_2_right_buffer_ccd_side_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_escape_err_signal                : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_escape_err_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_escape_err_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_indicate_signal               : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_rmap_target_indicate_o -> rmap_mem_ffee_deb_area:channel_hk_2_rmap_target_indicate_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_running_signal                   : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_running_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_running_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_credit_err_signal                : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_credit_err_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_credit_err_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_side_signal               : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_left_buffer_ccd_side_o -> rmap_mem_ffee_deb_area:channel_hk_2_left_buffer_ccd_side_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_err_right_buffer_overflow_signal          : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_err_right_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_2_err_right_buffer_overflow_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_status_signal                 : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:channel_hk_rmap_target_status_o -> rmap_mem_ffee_deb_area:channel_hk_2_rmap_target_status_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_parity_err_signal                : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_parity_err_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_parity_err_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_disconnect_signal                : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_disconnect_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_disconnect_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_connecting_signal                : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_connecting_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_connecting_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_started_signal                   : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_spw_link_started_o -> rmap_mem_ffee_deb_area:channel_hk_2_spw_link_started_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_number_signal            : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch3:channel_hk_right_buffer_ccd_number_o -> rmap_mem_ffee_deb_area:channel_hk_2_right_buffer_ccd_number_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_frame_counter_signal                      : std_logic_vector(15 downto 0);  -- Communication_Module_v2_Ch3:channel_hk_frame_counter_o -> rmap_mem_ffee_deb_area:channel_hk_2_frame_counter_i
	signal communication_module_v2_ch3_conduit_end_channel_hk_out_err_left_buffer_overflow_signal           : std_logic;                      -- Communication_Module_v2_Ch3:channel_hk_err_left_buffer_overflow_o -> rmap_mem_ffee_deb_area:channel_hk_2_err_left_buffer_overflow_i
	signal communication_module_v2_ch1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal          : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch1:channel_win_mem_addr_offset_o -> rmap_mem_ffee_deb_area:channel_win_mem_addr_offset_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_1_write_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_1_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_1_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_1_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_1_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_1_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_1_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb1_fee_hk_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_1_writedata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_5_write_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_5_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_5_rd_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_5_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_5_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_5_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_5_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb1_fee_hk_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_5_writedata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_7_write_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_7_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_7_rd_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_7_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_7_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_7_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_7_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb1_fee_hk_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_7_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_0_write_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_0_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_0_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_0_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_0_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_0_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_0_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb1_rmap_target_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_0_writedata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_2_write_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_2_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_2_rd_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_2_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_2_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_2_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_2_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb1_rmap_target_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_2_writedata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_3_write_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_3_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_3_rd_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_3_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_3_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_3_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_3_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb2_fee_hk_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_3_writedata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_5_write_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_5_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_5_rd_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_5_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_5_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_5_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_5_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb2_fee_hk_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_5_writedata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_7_write_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_7_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_7_rd_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_7_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_7_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_7_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_7_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb2_fee_hk_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_7_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_0_write_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_0_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_0_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_0_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_0_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_0_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_0_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb2_rmap_target_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_0_writedata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_3_write_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_3_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_3_rd_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_3_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_3_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_3_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_3_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb3_fee_hk_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_3_writedata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_5_write_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_5_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_5_rd_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_5_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_5_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_5_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_5_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb3_fee_hk_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_5_writedata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_7_write_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_7_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_7_rd_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_7_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_7_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_7_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_7_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb3_fee_hk_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_7_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_0_write_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_0_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_0_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_0_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_0_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_0_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_0_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb3_rmap_target_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_0_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_1_write_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_1_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_1_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_1_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_1_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_1_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_1_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb4_fee_hk_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_1_writedata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_3_write_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_3_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_3_rd_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_3_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_3_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_3_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_3_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb4_fee_hk_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_3_writedata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_5_write_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_5_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_5_rd_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_5_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_5_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_5_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_5_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb4_fee_hk_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_5_writedata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_7_write_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_7_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_7_rd_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_7_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_7_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_7_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_7_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb4_fee_hk_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_7_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_write_signal                  : std_logic;                      -- Communication_Module_v2_Ch1:rmm_deb_fee_hk_write_o -> rmap_mem_ffee_deb_area:rms_rmap_1_write_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_1_readdata_o -> Communication_Module_v2_Ch1:rmm_deb_fee_hk_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_deb_fee_hk_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_1_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_deb_fee_hk_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_1_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_read_signal                   : std_logic;                      -- Communication_Module_v2_Ch1:rmm_deb_fee_hk_read_o -> rmap_mem_ffee_deb_area:rms_rmap_1_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_1_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_deb_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_1_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_deb_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal              : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_deb_fee_hk_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_1_writedata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_write_signal                  : std_logic;                      -- Communication_Module_v2_Ch2:rmm_deb_fee_hk_write_o -> rmap_mem_ffee_deb_area:rms_rmap_3_write_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_3_readdata_o -> Communication_Module_v2_Ch2:rmm_deb_fee_hk_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_deb_fee_hk_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_3_rd_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_deb_fee_hk_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_3_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_read_signal                   : std_logic;                      -- Communication_Module_v2_Ch2:rmm_deb_fee_hk_read_o -> rmap_mem_ffee_deb_area:rms_rmap_3_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_3_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_deb_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_3_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_deb_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal              : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_deb_fee_hk_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_3_writedata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_write_signal                  : std_logic;                      -- Communication_Module_v2_Ch3:rmm_deb_fee_hk_write_o -> rmap_mem_ffee_deb_area:rms_rmap_5_write_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_5_readdata_o -> Communication_Module_v2_Ch3:rmm_deb_fee_hk_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_deb_fee_hk_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_5_rd_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_deb_fee_hk_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_5_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_read_signal                   : std_logic;                      -- Communication_Module_v2_Ch3:rmm_deb_fee_hk_read_o -> rmap_mem_ffee_deb_area:rms_rmap_5_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_5_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_deb_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_5_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_deb_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal              : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_deb_fee_hk_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_5_writedata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_write_signal                  : std_logic;                      -- Communication_Module_v2_Ch4:rmm_deb_fee_hk_write_o -> rmap_mem_ffee_deb_area:rms_rmap_7_write_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_7_readdata_o -> Communication_Module_v2_Ch4:rmm_deb_fee_hk_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_deb_fee_hk_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_7_rd_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal             : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_deb_fee_hk_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_7_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_read_signal                   : std_logic;                      -- Communication_Module_v2_Ch4:rmm_deb_fee_hk_read_o -> rmap_mem_ffee_deb_area:rms_rmap_7_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_7_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_deb_fee_hk_wr_waitrequest_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_7_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_deb_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal              : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_deb_fee_hk_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_7_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_write_signal             : std_logic;                      -- Communication_Module_v2_Ch1:rmm_deb_rmap_target_write_o -> rmap_mem_ffee_deb_area:rms_rmap_0_write_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_0_readdata_o -> Communication_Module_v2_Ch1:rmm_deb_rmap_target_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_deb_rmap_target_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_0_rd_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_deb_rmap_target_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_0_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_read_signal              : std_logic;                      -- Communication_Module_v2_Ch1:rmm_deb_rmap_target_read_o -> rmap_mem_ffee_deb_area:rms_rmap_0_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_0_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_deb_rmap_target_wr_waitrequest_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_0_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_deb_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal         : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_deb_rmap_target_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_0_writedata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_0_write_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_0_rd_address_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_0_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_0_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_0_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_0_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_0_writedata_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_0_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb4_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_1_write_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_1_rd_address_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_1_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_1_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_1_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_1_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_wr_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_1_writedata_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_1_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb2_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_1_write_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_1_rd_address_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_1_readdata_o -> Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_readdata_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_1_wr_address_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_1_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_1_wr_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_wr_waitrequest_i
	signal communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_1_writedata_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_1_rd_waitrequest_o -> Communication_Module_v2_Ch1:rmm_aeb3_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_2_write_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_2_rd_address_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_2_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_2_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_2_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_2_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_2_writedata_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_2_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb2_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_2_write_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_2_rd_address_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_2_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_2_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_2_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_2_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_2_writedata_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_2_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb3_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_2_write_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_2_rd_address_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_2_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_2_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_2_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_2_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_2_writedata_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_2_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb4_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_write_signal             : std_logic;                      -- Communication_Module_v2_Ch2:rmm_deb_rmap_target_write_o -> rmap_mem_ffee_deb_area:rms_rmap_2_write_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_deb_rmap_target_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_2_rd_address_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_2_readdata_o -> Communication_Module_v2_Ch2:rmm_deb_rmap_target_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_deb_rmap_target_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_2_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_read_signal              : std_logic;                      -- Communication_Module_v2_Ch2:rmm_deb_rmap_target_read_o -> rmap_mem_ffee_deb_area:rms_rmap_2_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_2_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_deb_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal         : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_deb_rmap_target_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_2_writedata_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_2_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_deb_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal                 : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_3_write_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_3_rd_address_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_3_readdata_o -> Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_readdata_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal            : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_3_wr_address_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal                  : std_logic;                      -- Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_3_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_3_wr_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_wr_waitrequest_i
	signal communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal             : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_3_writedata_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_3_rd_waitrequest_o -> Communication_Module_v2_Ch2:rmm_aeb1_fee_hk_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_4_write_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_4_rd_address_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_4_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_4_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_4_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_4_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_4_writedata_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_4_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb1_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_4_write_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_4_rd_address_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_4_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_4_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_4_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_4_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_4_writedata_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_4_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb2_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_4_write_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_4_rd_address_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_4_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_4_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_4_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_4_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_4_writedata_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_4_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb3_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_4_write_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_4_rd_address_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_4_readdata_o -> Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_4_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_4_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_4_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_4_writedata_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_4_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_aeb4_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_write_signal             : std_logic;                      -- Communication_Module_v2_Ch3:rmm_deb_rmap_target_write_o -> rmap_mem_ffee_deb_area:rms_rmap_4_write_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_deb_rmap_target_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_4_rd_address_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_4_readdata_o -> Communication_Module_v2_Ch3:rmm_deb_rmap_target_readdata_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:rmm_deb_rmap_target_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_4_wr_address_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_read_signal              : std_logic;                      -- Communication_Module_v2_Ch3:rmm_deb_rmap_target_read_o -> rmap_mem_ffee_deb_area:rms_rmap_4_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_4_wr_waitrequest_o -> Communication_Module_v2_Ch3:rmm_deb_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal         : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:rmm_deb_rmap_target_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_4_writedata_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_4_rd_waitrequest_o -> Communication_Module_v2_Ch3:rmm_deb_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_write_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_6_write_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_6_rd_address_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_1_area:rms_rmap_6_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_6_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_read_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_6_read_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_6_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_writedata_o -> rmap_mem_ffee_aeb_1_area:rms_rmap_6_writedata_i
	signal rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_1_area:rms_rmap_6_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb1_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_write_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_6_write_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_6_rd_address_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_2_area:rms_rmap_6_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_6_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_read_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_6_read_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_6_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_writedata_o -> rmap_mem_ffee_aeb_2_area:rms_rmap_6_writedata_i
	signal rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_2_area:rms_rmap_6_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb2_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_write_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_6_write_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_6_rd_address_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_3_area:rms_rmap_6_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_6_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_read_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_6_read_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_6_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_writedata_o -> rmap_mem_ffee_aeb_3_area:rms_rmap_6_writedata_i
	signal rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_3_area:rms_rmap_6_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb3_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal            : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_write_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_6_write_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_rd_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_6_rd_address_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_readdata_signal                            : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_aeb_4_area:rms_rmap_6_readdata_o -> Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal       : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_wr_address_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_6_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal             : std_logic;                      -- Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_read_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_6_read_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_6_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal        : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_writedata_o -> rmap_mem_ffee_aeb_4_area:rms_rmap_6_writedata_i
	signal rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal                      : std_logic;                      -- rmap_mem_ffee_aeb_4_area:rms_rmap_6_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_aeb4_rmap_target_rd_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_write_signal             : std_logic;                      -- Communication_Module_v2_Ch4:rmm_deb_rmap_target_write_o -> rmap_mem_ffee_deb_area:rms_rmap_6_write_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_deb_rmap_target_rd_address_o -> rmap_mem_ffee_deb_area:rms_rmap_6_rd_address_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_readdata_signal                              : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:rms_rmap_6_readdata_o -> Communication_Module_v2_Ch4:rmm_deb_rmap_target_readdata_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal        : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:rmm_deb_rmap_target_wr_address_o -> rmap_mem_ffee_deb_area:rms_rmap_6_wr_address_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_read_signal              : std_logic;                      -- Communication_Module_v2_Ch4:rmm_deb_rmap_target_read_o -> rmap_mem_ffee_deb_area:rms_rmap_6_read_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_6_wr_waitrequest_o -> Communication_Module_v2_Ch4:rmm_deb_rmap_target_wr_waitrequest_i
	signal communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal         : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:rmm_deb_rmap_target_writedata_o -> rmap_mem_ffee_deb_area:rms_rmap_6_writedata_i
	signal rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal                        : std_logic;                      -- rmap_mem_ffee_deb_area:rms_rmap_6_rd_waitrequest_o -> Communication_Module_v2_Ch4:rmm_deb_rmap_target_rd_waitrequest_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Demux_Ch2:spw_data_rx_status_rxvalid_o -> Communication_Module_v2_Ch2:spw_data_rx_status_rxvalid_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Demux_Ch2:spw_errinj_ctrl_errinj_busy_o -> Communication_Module_v2_Ch2:spw_errinj_ctrl_errinj_busy_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch2:spw_errinj_ctrl_start_errinj_o -> SpaceWire_Demux_Ch2:spw_errinj_ctrl_start_errinj_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:spw_data_tx_command_txdata_o -> SpaceWire_Demux_Ch2:spw_data_tx_command_txdata_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_error_errdisc_o -> Communication_Module_v2_Ch2:spw_link_error_errdisc_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch2:spw_data_tx_status_txhalff_o -> Communication_Module_v2_Ch2:spw_data_tx_status_txhalff_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  : std_logic;                      -- Communication_Module_v2_Ch2:spw_data_tx_command_txwrite_o -> SpaceWire_Demux_Ch2:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Demux_Ch2:spw_timecode_rx_tick_out_o -> Communication_Module_v2_Ch2:spw_timecode_rx_tick_out_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch2:spw_data_rx_status_rxhalff_o -> Communication_Module_v2_Ch2:spw_data_rx_status_rxhalff_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  : std_logic_vector(3 downto 0);   -- Communication_Module_v2_Ch2:spw_errinj_ctrl_errinj_code_o -> SpaceWire_Demux_Ch2:spw_errinj_ctrl_errinj_code_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch2:spw_timecode_rx_time_out_o -> Communication_Module_v2_Ch2:spw_timecode_rx_time_out_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_status_connecting_o -> Communication_Module_v2_Ch2:spw_link_status_connecting_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch2:spw_data_rx_status_rxdata_o -> Communication_Module_v2_Ch2:spw_data_rx_status_rxdata_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch2:spw_timecode_rx_ctrl_out_o -> Communication_Module_v2_Ch2:spw_timecode_rx_ctrl_out_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch2:spw_errinj_ctrl_reset_errinj_o -> SpaceWire_Demux_Ch2:spw_errinj_ctrl_reset_errinj_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   : std_logic;                      -- Communication_Module_v2_Ch2:spw_data_tx_command_txflag_o -> SpaceWire_Demux_Ch2:spw_data_tx_command_txflag_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   : std_logic;                      -- Communication_Module_v2_Ch2:spw_link_command_linkstart_o -> SpaceWire_Demux_Ch2:spw_link_command_linkstart_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   : std_logic;                      -- Communication_Module_v2_Ch2:spw_data_rx_command_rxread_o -> SpaceWire_Demux_Ch2:spw_data_rx_command_rxread_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_enable_signal      : std_logic;                      -- Communication_Module_v2_Ch2:spw_link_command_enable_o -> SpaceWire_Demux_Ch2:spw_link_command_enable_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_status_running_o -> Communication_Module_v2_Ch2:spw_link_status_running_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_status_started_o -> Communication_Module_v2_Ch2:spw_link_status_started_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_error_errpar_o -> Communication_Module_v2_Ch2:spw_link_error_errpar_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     : std_logic;                      -- Communication_Module_v2_Ch2:spw_link_command_linkdis_o -> SpaceWire_Demux_Ch2:spw_link_command_linkdis_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_error_erresc_o -> Communication_Module_v2_Ch2:spw_link_error_erresc_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Demux_Ch2:spw_data_tx_status_txrdy_o -> Communication_Module_v2_Ch2:spw_data_tx_status_txrdy_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      : std_logic;                      -- Communication_Module_v2_Ch2:spw_timecode_tx_tick_in_o -> SpaceWire_Demux_Ch2:spw_timecode_tx_tick_in_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch2:spw_link_command_txdivcnt_o -> SpaceWire_Demux_Ch2:spw_link_command_txdivcnt_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      : std_logic_vector(5 downto 0);   -- Communication_Module_v2_Ch2:spw_timecode_tx_time_in_o -> SpaceWire_Demux_Ch2:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Demux_Ch2:spw_data_rx_status_rxflag_o -> Communication_Module_v2_Ch2:spw_data_rx_status_rxflag_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch2:spw_timecode_tx_ctrl_in_o -> SpaceWire_Demux_Ch2:spw_timecode_tx_ctrl_in_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Demux_Ch2:spw_errinj_ctrl_errinj_ready_o -> Communication_Module_v2_Ch2:spw_errinj_ctrl_errinj_ready_i
	signal communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_autostart_signal   : std_logic;                      -- Communication_Module_v2_Ch2:spw_link_command_autostart_o -> SpaceWire_Demux_Ch2:spw_link_command_autostart_i
	signal spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Demux_Ch2:spw_link_error_errcred_o -> Communication_Module_v2_Ch2:spw_link_error_errcred_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_B:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch2:spw_ct0_data_rx_status_rxvalid_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_B:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch2:spw_ct0_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_B:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct0_data_tx_command_txdata_o -> SpaceWire_Channel_B:spw_data_tx_command_txdata_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_B:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch2:spw_ct0_link_error_errdisc_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_B:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch2:spw_ct0_data_tx_status_txhalff_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_data_tx_command_txwrite_o -> SpaceWire_Channel_B:spw_data_tx_command_txwrite_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_B:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch2:spw_ct0_timecode_rx_tick_out_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_B:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch2:spw_ct0_data_rx_status_rxhalff_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct0_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_B:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_B:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch2:spw_ct0_timecode_rx_time_out_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_B:spw_link_status_connecting_o -> SpaceWire_Demux_Ch2:spw_ct0_link_status_connecting_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_B:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch2:spw_ct0_data_rx_status_rxdata_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_B:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch2:spw_ct0_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_B:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_data_tx_command_txflag_o -> SpaceWire_Channel_B:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_link_command_linkstart_o -> SpaceWire_Channel_B:spw_link_command_linkstart_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_data_rx_command_rxread_o -> SpaceWire_Channel_B:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_link_command_enable_o -> SpaceWire_Channel_B:spw_link_command_enable_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_B:spw_link_status_running_o -> SpaceWire_Demux_Ch2:spw_ct0_link_status_running_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_B:spw_link_status_started_o -> SpaceWire_Demux_Ch2:spw_ct0_link_status_started_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_B:spw_link_error_errpar_o -> SpaceWire_Demux_Ch2:spw_ct0_link_error_errpar_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_link_command_linkdis_o -> SpaceWire_Channel_B:spw_link_command_linkdis_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_B:spw_link_error_erresc_o -> SpaceWire_Demux_Ch2:spw_ct0_link_error_erresc_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_B:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch2:spw_ct0_data_tx_status_txrdy_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_timecode_tx_tick_in_o -> SpaceWire_Channel_B:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct0_link_command_txdivcnt_o -> SpaceWire_Channel_B:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct0_timecode_tx_time_in_o -> SpaceWire_Channel_B:spw_timecode_tx_time_in_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_B:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch2:spw_ct0_data_rx_status_rxflag_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct0_timecode_tx_ctrl_in_o -> SpaceWire_Channel_B:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_B:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch2:spw_ct0_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct0_link_command_autostart_o -> SpaceWire_Channel_B:spw_link_command_autostart_i
	signal spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_B:spw_link_error_errcred_o -> SpaceWire_Demux_Ch2:spw_ct0_link_error_errcred_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_D:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch4:spw_ct0_data_rx_status_rxvalid_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_D:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch4:spw_ct0_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_D:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct0_data_tx_command_txdata_o -> SpaceWire_Channel_D:spw_data_tx_command_txdata_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_D:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch4:spw_ct0_link_error_errdisc_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_D:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch4:spw_ct0_data_tx_status_txhalff_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_data_tx_command_txwrite_o -> SpaceWire_Channel_D:spw_data_tx_command_txwrite_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_D:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch4:spw_ct0_timecode_rx_tick_out_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_D:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch4:spw_ct0_data_rx_status_rxhalff_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct0_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_D:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_D:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch4:spw_ct0_timecode_rx_time_out_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_D:spw_link_status_connecting_o -> SpaceWire_Demux_Ch4:spw_ct0_link_status_connecting_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_D:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch4:spw_ct0_data_rx_status_rxdata_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_D:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch4:spw_ct0_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_D:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_data_tx_command_txflag_o -> SpaceWire_Channel_D:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_link_command_linkstart_o -> SpaceWire_Channel_D:spw_link_command_linkstart_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_data_rx_command_rxread_o -> SpaceWire_Channel_D:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_link_command_enable_o -> SpaceWire_Channel_D:spw_link_command_enable_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_D:spw_link_status_running_o -> SpaceWire_Demux_Ch4:spw_ct0_link_status_running_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_D:spw_link_status_started_o -> SpaceWire_Demux_Ch4:spw_ct0_link_status_started_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_D:spw_link_error_errpar_o -> SpaceWire_Demux_Ch4:spw_ct0_link_error_errpar_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_link_command_linkdis_o -> SpaceWire_Channel_D:spw_link_command_linkdis_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_D:spw_link_error_erresc_o -> SpaceWire_Demux_Ch4:spw_ct0_link_error_erresc_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_D:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch4:spw_ct0_data_tx_status_txrdy_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_timecode_tx_tick_in_o -> SpaceWire_Channel_D:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct0_link_command_txdivcnt_o -> SpaceWire_Channel_D:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct0_timecode_tx_time_in_o -> SpaceWire_Channel_D:spw_timecode_tx_time_in_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_D:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch4:spw_ct0_data_rx_status_rxflag_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct0_timecode_tx_ctrl_in_o -> SpaceWire_Channel_D:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_D:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch4:spw_ct0_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct0_link_command_autostart_o -> SpaceWire_Channel_D:spw_link_command_autostart_i
	signal spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_D:spw_link_error_errcred_o -> SpaceWire_Demux_Ch4:spw_ct0_link_error_errcred_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_E:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch1:spw_ct1_data_rx_status_rxvalid_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_E:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch1:spw_ct1_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_E:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct1_data_tx_command_txdata_o -> SpaceWire_Channel_E:spw_data_tx_command_txdata_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_E:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch1:spw_ct1_link_error_errdisc_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_E:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch1:spw_ct1_data_tx_status_txhalff_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_data_tx_command_txwrite_o -> SpaceWire_Channel_E:spw_data_tx_command_txwrite_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_E:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch1:spw_ct1_timecode_rx_tick_out_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_E:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch1:spw_ct1_data_rx_status_rxhalff_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct1_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_E:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_E:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch1:spw_ct1_timecode_rx_time_out_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_E:spw_link_status_connecting_o -> SpaceWire_Demux_Ch1:spw_ct1_link_status_connecting_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_E:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch1:spw_ct1_data_rx_status_rxdata_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_E:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch1:spw_ct1_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_E:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_data_tx_command_txflag_o -> SpaceWire_Channel_E:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_link_command_linkstart_o -> SpaceWire_Channel_E:spw_link_command_linkstart_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_data_rx_command_rxread_o -> SpaceWire_Channel_E:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_link_command_enable_o -> SpaceWire_Channel_E:spw_link_command_enable_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_E:spw_link_status_running_o -> SpaceWire_Demux_Ch1:spw_ct1_link_status_running_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_E:spw_link_status_started_o -> SpaceWire_Demux_Ch1:spw_ct1_link_status_started_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_E:spw_link_error_errpar_o -> SpaceWire_Demux_Ch1:spw_ct1_link_error_errpar_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_link_command_linkdis_o -> SpaceWire_Channel_E:spw_link_command_linkdis_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_E:spw_link_error_erresc_o -> SpaceWire_Demux_Ch1:spw_ct1_link_error_erresc_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_E:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch1:spw_ct1_data_tx_status_txrdy_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_timecode_tx_tick_in_o -> SpaceWire_Channel_E:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct1_link_command_txdivcnt_o -> SpaceWire_Channel_E:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct1_timecode_tx_time_in_o -> SpaceWire_Channel_E:spw_timecode_tx_time_in_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_E:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch1:spw_ct1_data_rx_status_rxflag_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct1_timecode_tx_ctrl_in_o -> SpaceWire_Channel_E:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_E:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch1:spw_ct1_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct1_link_command_autostart_o -> SpaceWire_Channel_E:spw_link_command_autostart_i
	signal spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_E:spw_link_error_errcred_o -> SpaceWire_Demux_Ch1:spw_ct1_link_error_errcred_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Demux_Ch1:spw_data_rx_status_rxvalid_o -> Communication_Module_v2_Ch1:spw_data_rx_status_rxvalid_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Demux_Ch1:spw_errinj_ctrl_errinj_busy_o -> Communication_Module_v2_Ch1:spw_errinj_ctrl_errinj_busy_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch1:spw_errinj_ctrl_start_errinj_o -> SpaceWire_Demux_Ch1:spw_errinj_ctrl_start_errinj_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:spw_data_tx_command_txdata_o -> SpaceWire_Demux_Ch1:spw_data_tx_command_txdata_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_error_errdisc_o -> Communication_Module_v2_Ch1:spw_link_error_errdisc_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch1:spw_data_tx_status_txhalff_o -> Communication_Module_v2_Ch1:spw_data_tx_status_txhalff_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Demux_Ch1:spw_timecode_rx_tick_out_o -> Communication_Module_v2_Ch1:spw_timecode_rx_tick_out_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch1:spw_data_rx_status_rxhalff_o -> Communication_Module_v2_Ch1:spw_data_rx_status_rxhalff_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  : std_logic;                      -- Communication_Module_v2_Ch1:spw_data_tx_command_txwrite_o -> SpaceWire_Demux_Ch1:spw_data_tx_command_txwrite_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  : std_logic_vector(3 downto 0);   -- Communication_Module_v2_Ch1:spw_errinj_ctrl_errinj_code_o -> SpaceWire_Demux_Ch1:spw_errinj_ctrl_errinj_code_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch1:spw_timecode_rx_time_out_o -> Communication_Module_v2_Ch1:spw_timecode_rx_time_out_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_status_connecting_o -> Communication_Module_v2_Ch1:spw_link_status_connecting_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch1:spw_data_rx_status_rxdata_o -> Communication_Module_v2_Ch1:spw_data_rx_status_rxdata_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch1:spw_timecode_rx_ctrl_out_o -> Communication_Module_v2_Ch1:spw_timecode_rx_ctrl_out_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch1:spw_errinj_ctrl_reset_errinj_o -> SpaceWire_Demux_Ch1:spw_errinj_ctrl_reset_errinj_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   : std_logic;                      -- Communication_Module_v2_Ch1:spw_data_tx_command_txflag_o -> SpaceWire_Demux_Ch1:spw_data_tx_command_txflag_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   : std_logic;                      -- Communication_Module_v2_Ch1:spw_link_command_linkstart_o -> SpaceWire_Demux_Ch1:spw_link_command_linkstart_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   : std_logic;                      -- Communication_Module_v2_Ch1:spw_data_rx_command_rxread_o -> SpaceWire_Demux_Ch1:spw_data_rx_command_rxread_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_enable_signal      : std_logic;                      -- Communication_Module_v2_Ch1:spw_link_command_enable_o -> SpaceWire_Demux_Ch1:spw_link_command_enable_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_status_running_o -> Communication_Module_v2_Ch1:spw_link_status_running_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_status_started_o -> Communication_Module_v2_Ch1:spw_link_status_started_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_error_errpar_o -> Communication_Module_v2_Ch1:spw_link_error_errpar_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     : std_logic;                      -- Communication_Module_v2_Ch1:spw_link_command_linkdis_o -> SpaceWire_Demux_Ch1:spw_link_command_linkdis_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_error_erresc_o -> Communication_Module_v2_Ch1:spw_link_error_erresc_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Demux_Ch1:spw_data_tx_status_txrdy_o -> Communication_Module_v2_Ch1:spw_data_tx_status_txrdy_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      : std_logic;                      -- Communication_Module_v2_Ch1:spw_timecode_tx_tick_in_o -> SpaceWire_Demux_Ch1:spw_timecode_tx_tick_in_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch1:spw_link_command_txdivcnt_o -> SpaceWire_Demux_Ch1:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Demux_Ch1:spw_data_rx_status_rxflag_o -> Communication_Module_v2_Ch1:spw_data_rx_status_rxflag_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      : std_logic_vector(5 downto 0);   -- Communication_Module_v2_Ch1:spw_timecode_tx_time_in_o -> SpaceWire_Demux_Ch1:spw_timecode_tx_time_in_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch1:spw_timecode_tx_ctrl_in_o -> SpaceWire_Demux_Ch1:spw_timecode_tx_ctrl_in_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Demux_Ch1:spw_errinj_ctrl_errinj_ready_o -> Communication_Module_v2_Ch1:spw_errinj_ctrl_errinj_ready_i
	signal communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_autostart_signal   : std_logic;                      -- Communication_Module_v2_Ch1:spw_link_command_autostart_o -> SpaceWire_Demux_Ch1:spw_link_command_autostart_i
	signal spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Demux_Ch1:spw_link_error_errcred_o -> Communication_Module_v2_Ch1:spw_link_error_errcred_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Demux_Ch3:spw_data_rx_status_rxvalid_o -> Communication_Module_v2_Ch3:spw_data_rx_status_rxvalid_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Demux_Ch3:spw_errinj_ctrl_errinj_busy_o -> Communication_Module_v2_Ch3:spw_errinj_ctrl_errinj_busy_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch3:spw_errinj_ctrl_start_errinj_o -> SpaceWire_Demux_Ch3:spw_errinj_ctrl_start_errinj_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:spw_data_tx_command_txdata_o -> SpaceWire_Demux_Ch3:spw_data_tx_command_txdata_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_error_errdisc_o -> Communication_Module_v2_Ch3:spw_link_error_errdisc_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch3:spw_data_tx_status_txhalff_o -> Communication_Module_v2_Ch3:spw_data_tx_status_txhalff_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Demux_Ch3:spw_timecode_rx_tick_out_o -> Communication_Module_v2_Ch3:spw_timecode_rx_tick_out_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch3:spw_data_rx_status_rxhalff_o -> Communication_Module_v2_Ch3:spw_data_rx_status_rxhalff_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  : std_logic;                      -- Communication_Module_v2_Ch3:spw_data_tx_command_txwrite_o -> SpaceWire_Demux_Ch3:spw_data_tx_command_txwrite_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  : std_logic_vector(3 downto 0);   -- Communication_Module_v2_Ch3:spw_errinj_ctrl_errinj_code_o -> SpaceWire_Demux_Ch3:spw_errinj_ctrl_errinj_code_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch3:spw_timecode_rx_time_out_o -> Communication_Module_v2_Ch3:spw_timecode_rx_time_out_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_status_connecting_o -> Communication_Module_v2_Ch3:spw_link_status_connecting_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch3:spw_data_rx_status_rxdata_o -> Communication_Module_v2_Ch3:spw_data_rx_status_rxdata_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch3:spw_timecode_rx_ctrl_out_o -> Communication_Module_v2_Ch3:spw_timecode_rx_ctrl_out_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch3:spw_errinj_ctrl_reset_errinj_o -> SpaceWire_Demux_Ch3:spw_errinj_ctrl_reset_errinj_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   : std_logic;                      -- Communication_Module_v2_Ch3:spw_data_tx_command_txflag_o -> SpaceWire_Demux_Ch3:spw_data_tx_command_txflag_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   : std_logic;                      -- Communication_Module_v2_Ch3:spw_link_command_linkstart_o -> SpaceWire_Demux_Ch3:spw_link_command_linkstart_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   : std_logic;                      -- Communication_Module_v2_Ch3:spw_data_rx_command_rxread_o -> SpaceWire_Demux_Ch3:spw_data_rx_command_rxread_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_enable_signal      : std_logic;                      -- Communication_Module_v2_Ch3:spw_link_command_enable_o -> SpaceWire_Demux_Ch3:spw_link_command_enable_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_status_running_o -> Communication_Module_v2_Ch3:spw_link_status_running_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_status_started_o -> Communication_Module_v2_Ch3:spw_link_status_started_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_error_errpar_o -> Communication_Module_v2_Ch3:spw_link_error_errpar_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     : std_logic;                      -- Communication_Module_v2_Ch3:spw_link_command_linkdis_o -> SpaceWire_Demux_Ch3:spw_link_command_linkdis_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_error_erresc_o -> Communication_Module_v2_Ch3:spw_link_error_erresc_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Demux_Ch3:spw_data_tx_status_txrdy_o -> Communication_Module_v2_Ch3:spw_data_tx_status_txrdy_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      : std_logic;                      -- Communication_Module_v2_Ch3:spw_timecode_tx_tick_in_o -> SpaceWire_Demux_Ch3:spw_timecode_tx_tick_in_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch3:spw_link_command_txdivcnt_o -> SpaceWire_Demux_Ch3:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Demux_Ch3:spw_data_rx_status_rxflag_o -> Communication_Module_v2_Ch3:spw_data_rx_status_rxflag_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      : std_logic_vector(5 downto 0);   -- Communication_Module_v2_Ch3:spw_timecode_tx_time_in_o -> SpaceWire_Demux_Ch3:spw_timecode_tx_time_in_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch3:spw_timecode_tx_ctrl_in_o -> SpaceWire_Demux_Ch3:spw_timecode_tx_ctrl_in_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Demux_Ch3:spw_errinj_ctrl_errinj_ready_o -> Communication_Module_v2_Ch3:spw_errinj_ctrl_errinj_ready_i
	signal communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_autostart_signal   : std_logic;                      -- Communication_Module_v2_Ch3:spw_link_command_autostart_o -> SpaceWire_Demux_Ch3:spw_link_command_autostart_i
	signal spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Demux_Ch3:spw_link_error_errcred_o -> Communication_Module_v2_Ch3:spw_link_error_errcred_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Demux_Ch4:spw_data_rx_status_rxvalid_o -> Communication_Module_v2_Ch4:spw_data_rx_status_rxvalid_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Demux_Ch4:spw_errinj_ctrl_errinj_busy_o -> Communication_Module_v2_Ch4:spw_errinj_ctrl_errinj_busy_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch4:spw_errinj_ctrl_start_errinj_o -> SpaceWire_Demux_Ch4:spw_errinj_ctrl_start_errinj_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal   : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:spw_data_tx_command_txdata_o -> SpaceWire_Demux_Ch4:spw_data_tx_command_txdata_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_error_errdisc_o -> Communication_Module_v2_Ch4:spw_link_error_errdisc_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch4:spw_data_tx_status_txhalff_o -> Communication_Module_v2_Ch4:spw_data_tx_status_txhalff_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Demux_Ch4:spw_timecode_rx_tick_out_o -> Communication_Module_v2_Ch4:spw_timecode_rx_tick_out_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Demux_Ch4:spw_data_rx_status_rxhalff_o -> Communication_Module_v2_Ch4:spw_data_rx_status_rxhalff_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal  : std_logic;                      -- Communication_Module_v2_Ch4:spw_data_tx_command_txwrite_o -> SpaceWire_Demux_Ch4:spw_data_tx_command_txwrite_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal  : std_logic_vector(3 downto 0);   -- Communication_Module_v2_Ch4:spw_errinj_ctrl_errinj_code_o -> SpaceWire_Demux_Ch4:spw_errinj_ctrl_errinj_code_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch4:spw_timecode_rx_time_out_o -> Communication_Module_v2_Ch4:spw_timecode_rx_time_out_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_status_connecting_o -> Communication_Module_v2_Ch4:spw_link_status_connecting_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch4:spw_data_rx_status_rxdata_o -> Communication_Module_v2_Ch4:spw_data_rx_status_rxdata_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch4:spw_timecode_rx_ctrl_out_o -> Communication_Module_v2_Ch4:spw_timecode_rx_ctrl_out_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal : std_logic;                      -- Communication_Module_v2_Ch4:spw_errinj_ctrl_reset_errinj_o -> SpaceWire_Demux_Ch4:spw_errinj_ctrl_reset_errinj_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal   : std_logic;                      -- Communication_Module_v2_Ch4:spw_data_tx_command_txflag_o -> SpaceWire_Demux_Ch4:spw_data_tx_command_txflag_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal   : std_logic;                      -- Communication_Module_v2_Ch4:spw_link_command_linkstart_o -> SpaceWire_Demux_Ch4:spw_link_command_linkstart_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal   : std_logic;                      -- Communication_Module_v2_Ch4:spw_data_rx_command_rxread_o -> SpaceWire_Demux_Ch4:spw_data_rx_command_rxread_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_enable_signal      : std_logic;                      -- Communication_Module_v2_Ch4:spw_link_command_enable_o -> SpaceWire_Demux_Ch4:spw_link_command_enable_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_status_running_o -> Communication_Module_v2_Ch4:spw_link_status_running_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_status_started_o -> Communication_Module_v2_Ch4:spw_link_status_started_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_error_errpar_o -> Communication_Module_v2_Ch4:spw_link_error_errpar_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal     : std_logic;                      -- Communication_Module_v2_Ch4:spw_link_command_linkdis_o -> SpaceWire_Demux_Ch4:spw_link_command_linkdis_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_error_erresc_o -> Communication_Module_v2_Ch4:spw_link_error_erresc_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Demux_Ch4:spw_data_tx_status_txrdy_o -> Communication_Module_v2_Ch4:spw_data_tx_status_txrdy_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal      : std_logic;                      -- Communication_Module_v2_Ch4:spw_timecode_tx_tick_in_o -> SpaceWire_Demux_Ch4:spw_timecode_tx_tick_in_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal    : std_logic_vector(7 downto 0);   -- Communication_Module_v2_Ch4:spw_link_command_txdivcnt_o -> SpaceWire_Demux_Ch4:spw_link_command_txdivcnt_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Demux_Ch4:spw_data_rx_status_rxflag_o -> Communication_Module_v2_Ch4:spw_data_rx_status_rxflag_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal      : std_logic_vector(5 downto 0);   -- Communication_Module_v2_Ch4:spw_timecode_tx_time_in_o -> SpaceWire_Demux_Ch4:spw_timecode_tx_time_in_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal      : std_logic_vector(1 downto 0);   -- Communication_Module_v2_Ch4:spw_timecode_tx_ctrl_in_o -> SpaceWire_Demux_Ch4:spw_timecode_tx_ctrl_in_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Demux_Ch4:spw_errinj_ctrl_errinj_ready_o -> Communication_Module_v2_Ch4:spw_errinj_ctrl_errinj_ready_i
	signal communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_autostart_signal   : std_logic;                      -- Communication_Module_v2_Ch4:spw_link_command_autostart_o -> SpaceWire_Demux_Ch4:spw_link_command_autostart_i
	signal spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Demux_Ch4:spw_link_error_errcred_o -> Communication_Module_v2_Ch4:spw_link_error_errcred_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_A:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch1:spw_ct0_data_rx_status_rxvalid_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_A:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch1:spw_ct0_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_A:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct0_data_tx_command_txdata_o -> SpaceWire_Channel_A:spw_data_tx_command_txdata_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_A:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch1:spw_ct0_link_error_errdisc_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_A:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch1:spw_ct0_data_tx_status_txhalff_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_A:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch1:spw_ct0_timecode_rx_tick_out_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_A:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch1:spw_ct0_data_rx_status_rxhalff_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_data_tx_command_txwrite_o -> SpaceWire_Channel_A:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct0_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_A:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_A:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch1:spw_ct0_timecode_rx_time_out_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_A:spw_link_status_connecting_o -> SpaceWire_Demux_Ch1:spw_ct0_link_status_connecting_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_A:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch1:spw_ct0_data_rx_status_rxdata_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_A:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch1:spw_ct0_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_A:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_data_tx_command_txflag_o -> SpaceWire_Channel_A:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_link_command_linkstart_o -> SpaceWire_Channel_A:spw_link_command_linkstart_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_data_rx_command_rxread_o -> SpaceWire_Channel_A:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_link_command_enable_o -> SpaceWire_Channel_A:spw_link_command_enable_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_A:spw_link_status_running_o -> SpaceWire_Demux_Ch1:spw_ct0_link_status_running_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_A:spw_link_status_started_o -> SpaceWire_Demux_Ch1:spw_ct0_link_status_started_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_A:spw_link_error_errpar_o -> SpaceWire_Demux_Ch1:spw_ct0_link_error_errpar_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_link_command_linkdis_o -> SpaceWire_Channel_A:spw_link_command_linkdis_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_A:spw_link_error_erresc_o -> SpaceWire_Demux_Ch1:spw_ct0_link_error_erresc_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_A:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch1:spw_ct0_data_tx_status_txrdy_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_timecode_tx_tick_in_o -> SpaceWire_Channel_A:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct0_link_command_txdivcnt_o -> SpaceWire_Channel_A:spw_link_command_txdivcnt_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_A:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch1:spw_ct0_data_rx_status_rxflag_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct0_timecode_tx_time_in_o -> SpaceWire_Channel_A:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch1:spw_ct0_timecode_tx_ctrl_in_o -> SpaceWire_Channel_A:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_A:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch1:spw_ct0_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch1:spw_ct0_link_command_autostart_o -> SpaceWire_Channel_A:spw_link_command_autostart_i
	signal spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_A:spw_link_error_errcred_o -> SpaceWire_Demux_Ch1:spw_ct0_link_error_errcred_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_C:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch3:spw_ct0_data_rx_status_rxvalid_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_C:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch3:spw_ct0_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_C:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct0_data_tx_command_txdata_o -> SpaceWire_Channel_C:spw_data_tx_command_txdata_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_C:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch3:spw_ct0_link_error_errdisc_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_C:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch3:spw_ct0_data_tx_status_txhalff_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_C:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch3:spw_ct0_timecode_rx_tick_out_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_C:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch3:spw_ct0_data_rx_status_rxhalff_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_data_tx_command_txwrite_o -> SpaceWire_Channel_C:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct0_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_C:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_C:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch3:spw_ct0_timecode_rx_time_out_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_C:spw_link_status_connecting_o -> SpaceWire_Demux_Ch3:spw_ct0_link_status_connecting_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_C:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch3:spw_ct0_data_rx_status_rxdata_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_C:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch3:spw_ct0_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_C:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_data_tx_command_txflag_o -> SpaceWire_Channel_C:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_link_command_linkstart_o -> SpaceWire_Channel_C:spw_link_command_linkstart_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_data_rx_command_rxread_o -> SpaceWire_Channel_C:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_link_command_enable_o -> SpaceWire_Channel_C:spw_link_command_enable_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_C:spw_link_status_running_o -> SpaceWire_Demux_Ch3:spw_ct0_link_status_running_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_C:spw_link_status_started_o -> SpaceWire_Demux_Ch3:spw_ct0_link_status_started_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_C:spw_link_error_errpar_o -> SpaceWire_Demux_Ch3:spw_ct0_link_error_errpar_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_link_command_linkdis_o -> SpaceWire_Channel_C:spw_link_command_linkdis_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_C:spw_link_error_erresc_o -> SpaceWire_Demux_Ch3:spw_ct0_link_error_erresc_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_C:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch3:spw_ct0_data_tx_status_txrdy_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_timecode_tx_tick_in_o -> SpaceWire_Channel_C:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct0_link_command_txdivcnt_o -> SpaceWire_Channel_C:spw_link_command_txdivcnt_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_C:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch3:spw_ct0_data_rx_status_rxflag_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct0_timecode_tx_time_in_o -> SpaceWire_Channel_C:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct0_timecode_tx_ctrl_in_o -> SpaceWire_Channel_C:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_C:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch3:spw_ct0_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct0_link_command_autostart_o -> SpaceWire_Channel_C:spw_link_command_autostart_i
	signal spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_C:spw_link_error_errcred_o -> SpaceWire_Demux_Ch3:spw_ct0_link_error_errcred_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_F:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch2:spw_ct1_data_rx_status_rxvalid_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_F:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch2:spw_ct1_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_F:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct1_data_tx_command_txdata_o -> SpaceWire_Channel_F:spw_data_tx_command_txdata_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_F:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch2:spw_ct1_link_error_errdisc_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_F:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch2:spw_ct1_data_tx_status_txhalff_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_F:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch2:spw_ct1_timecode_rx_tick_out_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_F:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch2:spw_ct1_data_rx_status_rxhalff_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_data_tx_command_txwrite_o -> SpaceWire_Channel_F:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct1_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_F:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_F:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch2:spw_ct1_timecode_rx_time_out_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_F:spw_link_status_connecting_o -> SpaceWire_Demux_Ch2:spw_ct1_link_status_connecting_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_F:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch2:spw_ct1_data_rx_status_rxdata_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_F:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch2:spw_ct1_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_F:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_data_tx_command_txflag_o -> SpaceWire_Channel_F:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_link_command_linkstart_o -> SpaceWire_Channel_F:spw_link_command_linkstart_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_data_rx_command_rxread_o -> SpaceWire_Channel_F:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_link_command_enable_o -> SpaceWire_Channel_F:spw_link_command_enable_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_F:spw_link_status_running_o -> SpaceWire_Demux_Ch2:spw_ct1_link_status_running_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_F:spw_link_status_started_o -> SpaceWire_Demux_Ch2:spw_ct1_link_status_started_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_F:spw_link_error_errpar_o -> SpaceWire_Demux_Ch2:spw_ct1_link_error_errpar_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_link_command_linkdis_o -> SpaceWire_Channel_F:spw_link_command_linkdis_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_F:spw_link_error_erresc_o -> SpaceWire_Demux_Ch2:spw_ct1_link_error_erresc_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_F:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch2:spw_ct1_data_tx_status_txrdy_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_timecode_tx_tick_in_o -> SpaceWire_Channel_F:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct1_link_command_txdivcnt_o -> SpaceWire_Channel_F:spw_link_command_txdivcnt_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_F:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch2:spw_ct1_data_rx_status_rxflag_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct1_timecode_tx_time_in_o -> SpaceWire_Channel_F:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch2:spw_ct1_timecode_tx_ctrl_in_o -> SpaceWire_Channel_F:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_F:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch2:spw_ct1_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch2:spw_ct1_link_command_autostart_o -> SpaceWire_Channel_F:spw_link_command_autostart_i
	signal spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_F:spw_link_error_errcred_o -> SpaceWire_Demux_Ch2:spw_ct1_link_error_errcred_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_G:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch3:spw_ct1_data_rx_status_rxvalid_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_G:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch3:spw_ct1_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_G:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct1_data_tx_command_txdata_o -> SpaceWire_Channel_G:spw_data_tx_command_txdata_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_G:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch3:spw_ct1_link_error_errdisc_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_G:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch3:spw_ct1_data_tx_status_txhalff_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_G:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch3:spw_ct1_timecode_rx_tick_out_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_G:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch3:spw_ct1_data_rx_status_rxhalff_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_data_tx_command_txwrite_o -> SpaceWire_Channel_G:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct1_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_G:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_G:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch3:spw_ct1_timecode_rx_time_out_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_G:spw_link_status_connecting_o -> SpaceWire_Demux_Ch3:spw_ct1_link_status_connecting_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_G:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch3:spw_ct1_data_rx_status_rxdata_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_G:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch3:spw_ct1_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_G:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_data_tx_command_txflag_o -> SpaceWire_Channel_G:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_link_command_linkstart_o -> SpaceWire_Channel_G:spw_link_command_linkstart_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_data_rx_command_rxread_o -> SpaceWire_Channel_G:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_link_command_enable_o -> SpaceWire_Channel_G:spw_link_command_enable_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_G:spw_link_status_running_o -> SpaceWire_Demux_Ch3:spw_ct1_link_status_running_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_G:spw_link_status_started_o -> SpaceWire_Demux_Ch3:spw_ct1_link_status_started_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_G:spw_link_error_errpar_o -> SpaceWire_Demux_Ch3:spw_ct1_link_error_errpar_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_link_command_linkdis_o -> SpaceWire_Channel_G:spw_link_command_linkdis_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_G:spw_link_error_erresc_o -> SpaceWire_Demux_Ch3:spw_ct1_link_error_erresc_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_G:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch3:spw_ct1_data_tx_status_txrdy_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_timecode_tx_tick_in_o -> SpaceWire_Channel_G:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct1_link_command_txdivcnt_o -> SpaceWire_Channel_G:spw_link_command_txdivcnt_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_G:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch3:spw_ct1_data_rx_status_rxflag_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct1_timecode_tx_time_in_o -> SpaceWire_Channel_G:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch3:spw_ct1_timecode_tx_ctrl_in_o -> SpaceWire_Channel_G:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_G:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch3:spw_ct1_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch3:spw_ct1_link_command_autostart_o -> SpaceWire_Channel_G:spw_link_command_autostart_i
	signal spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_G:spw_link_error_errcred_o -> SpaceWire_Demux_Ch3:spw_ct1_link_error_errcred_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal              : std_logic;                      -- SpaceWire_Channel_H:spw_data_rx_status_rxvalid_o -> SpaceWire_Demux_Ch4:spw_ct1_data_rx_status_rxvalid_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal             : std_logic;                      -- SpaceWire_Channel_H:spw_errinj_ctrl_errinj_busy_o -> SpaceWire_Demux_Ch4:spw_ct1_errinj_ctrl_errinj_busy_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_errinj_ctrl_start_errinj_o -> SpaceWire_Channel_H:spw_errinj_ctrl_start_errinj_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal         : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct1_data_tx_command_txdata_o -> SpaceWire_Channel_H:spw_data_tx_command_txdata_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal                  : std_logic;                      -- SpaceWire_Channel_H:spw_link_error_errdisc_o -> SpaceWire_Demux_Ch4:spw_ct1_link_error_errdisc_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal              : std_logic;                      -- SpaceWire_Channel_H:spw_data_tx_status_txhalff_o -> SpaceWire_Demux_Ch4:spw_ct1_data_tx_status_txhalff_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal                : std_logic;                      -- SpaceWire_Channel_H:spw_timecode_rx_tick_out_o -> SpaceWire_Demux_Ch4:spw_ct1_timecode_rx_tick_out_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal              : std_logic;                      -- SpaceWire_Channel_H:spw_data_rx_status_rxhalff_o -> SpaceWire_Demux_Ch4:spw_ct1_data_rx_status_rxhalff_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal        : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_data_tx_command_txwrite_o -> SpaceWire_Channel_H:spw_data_tx_command_txwrite_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal        : std_logic_vector(3 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct1_errinj_ctrl_errinj_code_o -> SpaceWire_Channel_H:spw_errinj_ctrl_errinj_code_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal                : std_logic_vector(5 downto 0);   -- SpaceWire_Channel_H:spw_timecode_rx_time_out_o -> SpaceWire_Demux_Ch4:spw_ct1_timecode_rx_time_out_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal              : std_logic;                      -- SpaceWire_Channel_H:spw_link_status_connecting_o -> SpaceWire_Demux_Ch4:spw_ct1_link_status_connecting_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal               : std_logic_vector(7 downto 0);   -- SpaceWire_Channel_H:spw_data_rx_status_rxdata_o -> SpaceWire_Demux_Ch4:spw_ct1_data_rx_status_rxdata_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal                : std_logic_vector(1 downto 0);   -- SpaceWire_Channel_H:spw_timecode_rx_ctrl_out_o -> SpaceWire_Demux_Ch4:spw_ct1_timecode_rx_ctrl_out_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal       : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_errinj_ctrl_reset_errinj_o -> SpaceWire_Channel_H:spw_errinj_ctrl_reset_errinj_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_data_tx_command_txflag_o -> SpaceWire_Channel_H:spw_data_tx_command_txflag_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_link_command_linkstart_o -> SpaceWire_Channel_H:spw_link_command_linkstart_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_data_rx_command_rxread_o -> SpaceWire_Channel_H:spw_data_rx_command_rxread_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_enable_signal            : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_link_command_enable_o -> SpaceWire_Channel_H:spw_link_command_enable_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal                 : std_logic;                      -- SpaceWire_Channel_H:spw_link_status_running_o -> SpaceWire_Demux_Ch4:spw_ct1_link_status_running_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal                 : std_logic;                      -- SpaceWire_Channel_H:spw_link_status_started_o -> SpaceWire_Demux_Ch4:spw_ct1_link_status_started_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal                   : std_logic;                      -- SpaceWire_Channel_H:spw_link_error_errpar_o -> SpaceWire_Demux_Ch4:spw_ct1_link_error_errpar_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal           : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_link_command_linkdis_o -> SpaceWire_Channel_H:spw_link_command_linkdis_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal                   : std_logic;                      -- SpaceWire_Channel_H:spw_link_error_erresc_o -> SpaceWire_Demux_Ch4:spw_ct1_link_error_erresc_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal                : std_logic;                      -- SpaceWire_Channel_H:spw_data_tx_status_txrdy_o -> SpaceWire_Demux_Ch4:spw_ct1_data_tx_status_txrdy_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal            : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_timecode_tx_tick_in_o -> SpaceWire_Channel_H:spw_timecode_tx_tick_in_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal          : std_logic_vector(7 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct1_link_command_txdivcnt_o -> SpaceWire_Channel_H:spw_link_command_txdivcnt_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal               : std_logic;                      -- SpaceWire_Channel_H:spw_data_rx_status_rxflag_o -> SpaceWire_Demux_Ch4:spw_ct1_data_rx_status_rxflag_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal            : std_logic_vector(5 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct1_timecode_tx_time_in_o -> SpaceWire_Channel_H:spw_timecode_tx_time_in_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal            : std_logic_vector(1 downto 0);   -- SpaceWire_Demux_Ch4:spw_ct1_timecode_tx_ctrl_in_o -> SpaceWire_Channel_H:spw_timecode_tx_ctrl_in_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal            : std_logic;                      -- SpaceWire_Channel_H:spw_errinj_ctrl_errinj_ready_o -> SpaceWire_Demux_Ch4:spw_ct1_errinj_ctrl_errinj_ready_i
	signal spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal         : std_logic;                      -- SpaceWire_Demux_Ch4:spw_ct1_link_command_autostart_o -> SpaceWire_Channel_H:spw_link_command_autostart_i
	signal spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal                  : std_logic;                      -- SpaceWire_Channel_H:spw_link_error_errcred_o -> SpaceWire_Demux_Ch4:spw_ct1_link_error_errcred_i
	signal ext_flash_tcm_data_outen                                                                         : std_logic;                      -- ext_flash:tcm_data_outen -> tristate_conduit_bridge_0:tcs_tcm_data_outen
	signal ext_flash_tcm_request                                                                            : std_logic;                      -- ext_flash:tcm_request -> tristate_conduit_bridge_0:request
	signal ext_flash_tcm_write_n_out                                                                        : std_logic;                      -- ext_flash:tcm_write_n_out -> tristate_conduit_bridge_0:tcs_tcm_write_n_out
	signal ext_flash_tcm_read_n_out                                                                         : std_logic;                      -- ext_flash:tcm_read_n_out -> tristate_conduit_bridge_0:tcs_tcm_read_n_out
	signal ext_flash_tcm_grant                                                                              : std_logic;                      -- tristate_conduit_bridge_0:grant -> ext_flash:tcm_grant
	signal ext_flash_tcm_chipselect_n_out                                                                   : std_logic;                      -- ext_flash:tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_tcm_chipselect_n_out
	signal ext_flash_tcm_address_out                                                                        : std_logic_vector(25 downto 0);  -- ext_flash:tcm_address_out -> tristate_conduit_bridge_0:tcs_tcm_address_out
	signal ext_flash_tcm_data_out                                                                           : std_logic_vector(15 downto 0);  -- ext_flash:tcm_data_out -> tristate_conduit_bridge_0:tcs_tcm_data_out
	signal ext_flash_tcm_data_in                                                                            : std_logic_vector(15 downto 0);  -- tristate_conduit_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	signal ftdi_umft601a_module_avalon_imgt_master_data_waitrequest                                         : std_logic;                      -- mm_interconnect_0:FTDI_UMFT601A_Module_avalon_imgt_master_data_waitrequest -> FTDI_UMFT601A_Module:avalon_imgt_master_data_waitrequest_i
	signal ftdi_umft601a_module_avalon_imgt_master_data_address                                             : std_logic_vector(63 downto 0);  -- FTDI_UMFT601A_Module:avalon_imgt_master_data_address_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_imgt_master_data_address
	signal ftdi_umft601a_module_avalon_imgt_master_data_write                                               : std_logic;                      -- FTDI_UMFT601A_Module:avalon_imgt_master_data_write_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_imgt_master_data_write
	signal ftdi_umft601a_module_avalon_imgt_master_data_writedata                                           : std_logic_vector(15 downto 0);  -- FTDI_UMFT601A_Module:avalon_imgt_master_data_writedata_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_imgt_master_data_writedata
	signal ftdi_umft601a_module_avalon_master_data_readdata                                                 : std_logic_vector(255 downto 0); -- mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_readdata -> FTDI_UMFT601A_Module:avalon_master_data_readdata_i
	signal ftdi_umft601a_module_avalon_master_data_waitrequest                                              : std_logic;                      -- mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_waitrequest -> FTDI_UMFT601A_Module:avalon_master_data_waitrequest_i
	signal ftdi_umft601a_module_avalon_master_data_address                                                  : std_logic_vector(63 downto 0);  -- FTDI_UMFT601A_Module:avalon_master_data_address_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_address
	signal ftdi_umft601a_module_avalon_master_data_read                                                     : std_logic;                      -- FTDI_UMFT601A_Module:avalon_master_data_read_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_read
	signal ftdi_umft601a_module_avalon_master_data_write                                                    : std_logic;                      -- FTDI_UMFT601A_Module:avalon_master_data_write_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_write
	signal ftdi_umft601a_module_avalon_master_data_writedata                                                : std_logic_vector(255 downto 0); -- FTDI_UMFT601A_Module:avalon_master_data_writedata_o -> mm_interconnect_0:FTDI_UMFT601A_Module_avalon_master_data_writedata
	signal memory_filler_avalon_master_data_waitrequest                                                     : std_logic;                      -- mm_interconnect_0:Memory_Filler_avalon_master_data_waitrequest -> Memory_Filler:avalon_master_data_waitrequest_i
	signal memory_filler_avalon_master_data_address                                                         : std_logic_vector(63 downto 0);  -- Memory_Filler:avalon_master_data_address_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_address
	signal memory_filler_avalon_master_data_write                                                           : std_logic;                      -- Memory_Filler:avalon_master_data_write_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_write
	signal memory_filler_avalon_master_data_writedata                                                       : std_logic_vector(255 downto 0); -- Memory_Filler:avalon_master_data_writedata_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_writedata
	signal communication_module_v2_ch1_avalon_mm_left_buffer_master_readdata                                : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_readdata -> Communication_Module_v2_Ch1:avm_left_buffer_readdata_i
	signal communication_module_v2_ch1_avalon_mm_left_buffer_master_waitrequest                             : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_waitrequest -> Communication_Module_v2_Ch1:avm_left_buffer_waitrequest_i
	signal communication_module_v2_ch1_avalon_mm_left_buffer_master_address                                 : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch1:avm_left_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_address
	signal communication_module_v2_ch1_avalon_mm_left_buffer_master_read                                    : std_logic;                      -- Communication_Module_v2_Ch1:avm_left_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_read
	signal communication_module_v2_ch2_avalon_mm_left_buffer_master_readdata                                : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_readdata -> Communication_Module_v2_Ch2:avm_left_buffer_readdata_i
	signal communication_module_v2_ch2_avalon_mm_left_buffer_master_waitrequest                             : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_waitrequest -> Communication_Module_v2_Ch2:avm_left_buffer_waitrequest_i
	signal communication_module_v2_ch2_avalon_mm_left_buffer_master_address                                 : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch2:avm_left_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_address
	signal communication_module_v2_ch2_avalon_mm_left_buffer_master_read                                    : std_logic;                      -- Communication_Module_v2_Ch2:avm_left_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_read
	signal communication_module_v2_ch4_avalon_mm_left_buffer_master_readdata                                : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_readdata -> Communication_Module_v2_Ch4:avm_left_buffer_readdata_i
	signal communication_module_v2_ch4_avalon_mm_left_buffer_master_waitrequest                             : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_waitrequest -> Communication_Module_v2_Ch4:avm_left_buffer_waitrequest_i
	signal communication_module_v2_ch4_avalon_mm_left_buffer_master_address                                 : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch4:avm_left_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_address
	signal communication_module_v2_ch4_avalon_mm_left_buffer_master_read                                    : std_logic;                      -- Communication_Module_v2_Ch4:avm_left_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_read
	signal communication_module_v2_ch3_avalon_mm_left_buffer_master_readdata                                : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_readdata -> Communication_Module_v2_Ch3:avm_left_buffer_readdata_i
	signal communication_module_v2_ch3_avalon_mm_left_buffer_master_waitrequest                             : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_waitrequest -> Communication_Module_v2_Ch3:avm_left_buffer_waitrequest_i
	signal communication_module_v2_ch3_avalon_mm_left_buffer_master_address                                 : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch3:avm_left_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_address
	signal communication_module_v2_ch3_avalon_mm_left_buffer_master_read                                    : std_logic;                      -- Communication_Module_v2_Ch3:avm_left_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_read
	signal communication_module_v2_ch1_avalon_mm_right_buffer_master_readdata                               : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_readdata -> Communication_Module_v2_Ch1:avm_right_buffer_readdata_i
	signal communication_module_v2_ch1_avalon_mm_right_buffer_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_waitrequest -> Communication_Module_v2_Ch1:avm_right_buffer_waitrequest_i
	signal communication_module_v2_ch1_avalon_mm_right_buffer_master_address                                : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch1:avm_right_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_address
	signal communication_module_v2_ch1_avalon_mm_right_buffer_master_read                                   : std_logic;                      -- Communication_Module_v2_Ch1:avm_right_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_read
	signal communication_module_v2_ch2_avalon_mm_right_buffer_master_readdata                               : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_readdata -> Communication_Module_v2_Ch2:avm_right_buffer_readdata_i
	signal communication_module_v2_ch2_avalon_mm_right_buffer_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_waitrequest -> Communication_Module_v2_Ch2:avm_right_buffer_waitrequest_i
	signal communication_module_v2_ch2_avalon_mm_right_buffer_master_address                                : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch2:avm_right_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_address
	signal communication_module_v2_ch2_avalon_mm_right_buffer_master_read                                   : std_logic;                      -- Communication_Module_v2_Ch2:avm_right_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_read
	signal communication_module_v2_ch4_avalon_mm_right_buffer_master_readdata                               : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_readdata -> Communication_Module_v2_Ch4:avm_right_buffer_readdata_i
	signal communication_module_v2_ch4_avalon_mm_right_buffer_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_waitrequest -> Communication_Module_v2_Ch4:avm_right_buffer_waitrequest_i
	signal communication_module_v2_ch4_avalon_mm_right_buffer_master_address                                : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch4:avm_right_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_address
	signal communication_module_v2_ch4_avalon_mm_right_buffer_master_read                                   : std_logic;                      -- Communication_Module_v2_Ch4:avm_right_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_read
	signal communication_module_v2_ch3_avalon_mm_right_buffer_master_readdata                               : std_logic_vector(255 downto 0); -- mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_readdata -> Communication_Module_v2_Ch3:avm_right_buffer_readdata_i
	signal communication_module_v2_ch3_avalon_mm_right_buffer_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_waitrequest -> Communication_Module_v2_Ch3:avm_right_buffer_waitrequest_i
	signal communication_module_v2_ch3_avalon_mm_right_buffer_master_address                                : std_logic_vector(63 downto 0);  -- Communication_Module_v2_Ch3:avm_right_buffer_address_o -> mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_address
	signal communication_module_v2_ch3_avalon_mm_right_buffer_master_read                                   : std_logic;                      -- Communication_Module_v2_Ch3:avm_right_buffer_read_o -> mm_interconnect_0:Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_read
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata                                            : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata -> rmap_mem_ffee_deb_area:avm_rmap_readdata_i
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest                                         : std_logic;                      -- mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest -> rmap_mem_ffee_deb_area:avm_rmap_waitrequest_i
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address                                             : std_logic_vector(63 downto 0);  -- rmap_mem_ffee_deb_area:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read                                                : std_logic;                      -- rmap_mem_ffee_deb_area:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write                                               : std_logic;                      -- rmap_mem_ffee_deb_area:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write
	signal rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata                                           : std_logic_vector(7 downto 0);   -- rmap_mem_ffee_deb_area:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata
	signal ddr2_address_span_extender_expanded_master_waitrequest                                           : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_waitrequest -> ddr2_address_span_extender:avm_m0_waitrequest
	signal ddr2_address_span_extender_expanded_master_readdata                                              : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdata -> ddr2_address_span_extender:avm_m0_readdata
	signal ddr2_address_span_extender_expanded_master_address                                               : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_address -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_address
	signal ddr2_address_span_extender_expanded_master_read                                                  : std_logic;                      -- ddr2_address_span_extender:avm_m0_read -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_read
	signal ddr2_address_span_extender_expanded_master_byteenable                                            : std_logic_vector(3 downto 0);   -- ddr2_address_span_extender:avm_m0_byteenable -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_byteenable
	signal ddr2_address_span_extender_expanded_master_readdatavalid                                         : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdatavalid -> ddr2_address_span_extender:avm_m0_readdatavalid
	signal ddr2_address_span_extender_expanded_master_write                                                 : std_logic;                      -- ddr2_address_span_extender:avm_m0_write -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_write
	signal ddr2_address_span_extender_expanded_master_writedata                                             : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_writedata -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_writedata
	signal ddr2_address_span_extender_expanded_master_burstcount                                            : std_logic_vector(7 downto 0);   -- ddr2_address_span_extender:avm_m0_burstcount -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_burstcount
	signal mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer                                          : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_beginbursttransfer -> m2_ddr2_memory:avl_burstbegin
	signal mm_interconnect_0_m2_ddr2_memory_avl_readdata                                                    : std_logic_vector(255 downto 0); -- m2_ddr2_memory:avl_rdata -> mm_interconnect_0:m2_ddr2_memory_avl_readdata
	signal m2_ddr2_memory_avl_waitrequest                                                                   : std_logic;                      -- m2_ddr2_memory:avl_ready -> m2_ddr2_memory_avl_waitrequest:in
	signal mm_interconnect_0_m2_ddr2_memory_avl_address                                                     : std_logic_vector(25 downto 0);  -- mm_interconnect_0:m2_ddr2_memory_avl_address -> m2_ddr2_memory:avl_addr
	signal mm_interconnect_0_m2_ddr2_memory_avl_read                                                        : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_read -> m2_ddr2_memory:avl_read_req
	signal mm_interconnect_0_m2_ddr2_memory_avl_byteenable                                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:m2_ddr2_memory_avl_byteenable -> m2_ddr2_memory:avl_be
	signal mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid                                               : std_logic;                      -- m2_ddr2_memory:avl_rdata_valid -> mm_interconnect_0:m2_ddr2_memory_avl_readdatavalid
	signal mm_interconnect_0_m2_ddr2_memory_avl_write                                                       : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_write -> m2_ddr2_memory:avl_write_req
	signal mm_interconnect_0_m2_ddr2_memory_avl_writedata                                                   : std_logic_vector(255 downto 0); -- mm_interconnect_0:m2_ddr2_memory_avl_writedata -> m2_ddr2_memory:avl_wdata
	signal mm_interconnect_0_m2_ddr2_memory_avl_burstcount                                                  : std_logic_vector(7 downto 0);   -- mm_interconnect_0:m2_ddr2_memory_avl_burstcount -> m2_ddr2_memory:avl_size
	signal mm_interconnect_0_m1_clock_bridge_s0_readdata                                                    : std_logic_vector(255 downto 0); -- m1_clock_bridge:s0_readdata -> mm_interconnect_0:m1_clock_bridge_s0_readdata
	signal mm_interconnect_0_m1_clock_bridge_s0_waitrequest                                                 : std_logic;                      -- m1_clock_bridge:s0_waitrequest -> mm_interconnect_0:m1_clock_bridge_s0_waitrequest
	signal mm_interconnect_0_m1_clock_bridge_s0_debugaccess                                                 : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_debugaccess -> m1_clock_bridge:s0_debugaccess
	signal mm_interconnect_0_m1_clock_bridge_s0_address                                                     : std_logic_vector(30 downto 0);  -- mm_interconnect_0:m1_clock_bridge_s0_address -> m1_clock_bridge:s0_address
	signal mm_interconnect_0_m1_clock_bridge_s0_read                                                        : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_read -> m1_clock_bridge:s0_read
	signal mm_interconnect_0_m1_clock_bridge_s0_byteenable                                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:m1_clock_bridge_s0_byteenable -> m1_clock_bridge:s0_byteenable
	signal mm_interconnect_0_m1_clock_bridge_s0_readdatavalid                                               : std_logic;                      -- m1_clock_bridge:s0_readdatavalid -> mm_interconnect_0:m1_clock_bridge_s0_readdatavalid
	signal mm_interconnect_0_m1_clock_bridge_s0_write                                                       : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_write -> m1_clock_bridge:s0_write
	signal mm_interconnect_0_m1_clock_bridge_s0_writedata                                                   : std_logic_vector(255 downto 0); -- mm_interconnect_0:m1_clock_bridge_s0_writedata -> m1_clock_bridge:s0_writedata
	signal mm_interconnect_0_m1_clock_bridge_s0_burstcount                                                  : std_logic_vector(2 downto 0);   -- mm_interconnect_0:m1_clock_bridge_s0_burstcount -> m1_clock_bridge:s0_burstcount
	signal nios2_gen2_0_data_master_readdata                                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                                             : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                                             : std_logic;                      -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                                 : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                                              : std_logic_vector(3 downto 0);   -- nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                                    : std_logic;                      -- nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                                   : std_logic;                      -- nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                                               : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                                      : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                                          : std_logic_vector(31 downto 0);  -- nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                                             : std_logic;                      -- nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                                                    : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal nios2_gen2_0_instruction_master_burstcount                                                       : std_logic_vector(3 downto 0);   -- nios2_gen2_0:i_burstcount -> mm_interconnect_1:nios2_gen2_0_instruction_master_burstcount
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect                                       : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata                                         : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest                                      : std_logic;                      -- jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address                                          : std_logic_vector(0 downto 0);   -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read                                             : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write                                            : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_readdata                    : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch1:avs_config_readdata_o -> mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_readdata
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_waitrequest                 : std_logic;                      -- Communication_Module_v2_Ch1:avs_config_waitrequest_o -> mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_waitrequest
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_address                     : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_address -> Communication_Module_v2_Ch1:avs_config_address_i
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_read                        : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_read -> Communication_Module_v2_Ch1:avs_config_read_i
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_write                       : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_write -> Communication_Module_v2_Ch1:avs_config_write_i
	signal mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Communication_Module_v2_Ch1_avalon_mm_config_slave_writedata -> Communication_Module_v2_Ch1:avs_config_writedata_i
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_readdata                    : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch2:avs_config_readdata_o -> mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_readdata
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_waitrequest                 : std_logic;                      -- Communication_Module_v2_Ch2:avs_config_waitrequest_o -> mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_waitrequest
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_address                     : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_address -> Communication_Module_v2_Ch2:avs_config_address_i
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_read                        : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_read -> Communication_Module_v2_Ch2:avs_config_read_i
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_write                       : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_write -> Communication_Module_v2_Ch2:avs_config_write_i
	signal mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Communication_Module_v2_Ch2_avalon_mm_config_slave_writedata -> Communication_Module_v2_Ch2:avs_config_writedata_i
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_readdata                    : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch4:avs_config_readdata_o -> mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_readdata
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_waitrequest                 : std_logic;                      -- Communication_Module_v2_Ch4:avs_config_waitrequest_o -> mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_waitrequest
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_address                     : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_address -> Communication_Module_v2_Ch4:avs_config_address_i
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_read                        : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_read -> Communication_Module_v2_Ch4:avs_config_read_i
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_write                       : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_write -> Communication_Module_v2_Ch4:avs_config_write_i
	signal mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Communication_Module_v2_Ch4_avalon_mm_config_slave_writedata -> Communication_Module_v2_Ch4:avs_config_writedata_i
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_readdata                    : std_logic_vector(31 downto 0);  -- Communication_Module_v2_Ch3:avs_config_readdata_o -> mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_readdata
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_waitrequest                 : std_logic;                      -- Communication_Module_v2_Ch3:avs_config_waitrequest_o -> mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_waitrequest
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_address                     : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_address -> Communication_Module_v2_Ch3:avs_config_address_i
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_read                        : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_read -> Communication_Module_v2_Ch3:avs_config_read_i
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_write                       : std_logic;                      -- mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_write -> Communication_Module_v2_Ch3:avs_config_write_i
	signal mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Communication_Module_v2_Ch3_avalon_mm_config_slave_writedata -> Communication_Module_v2_Ch3:avs_config_writedata_i
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata                            : std_logic_vector(31 downto 0);  -- rmap_mem_ffee_deb_area:avs_rmap_0_readdata_o -> mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest                         : std_logic;                      -- rmap_mem_ffee_deb_area:avs_rmap_0_waitrequest_o -> mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address                             : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address -> rmap_mem_ffee_deb_area:avs_rmap_0_address_i
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read                                : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read -> rmap_mem_ffee_deb_area:avs_rmap_0_read_i
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write                               : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write -> rmap_mem_ffee_deb_area:avs_rmap_0_write_i
	signal mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata                           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata -> rmap_mem_ffee_deb_area:avs_rmap_0_writedata_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata                          : std_logic_vector(31 downto 0);  -- rmap_mem_ffee_aeb_1_area:avs_rmap_0_readdata_o -> mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest                       : std_logic;                      -- rmap_mem_ffee_aeb_1_area:avs_rmap_0_waitrequest_o -> mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address -> rmap_mem_ffee_aeb_1_area:avs_rmap_0_address_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read                              : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read -> rmap_mem_ffee_aeb_1_area:avs_rmap_0_read_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write                             : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write -> rmap_mem_ffee_aeb_1_area:avs_rmap_0_write_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata -> rmap_mem_ffee_aeb_1_area:avs_rmap_0_writedata_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata                          : std_logic_vector(31 downto 0);  -- rmap_mem_ffee_aeb_2_area:avs_rmap_0_readdata_o -> mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest                       : std_logic;                      -- rmap_mem_ffee_aeb_2_area:avs_rmap_0_waitrequest_o -> mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address -> rmap_mem_ffee_aeb_2_area:avs_rmap_0_address_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read                              : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read -> rmap_mem_ffee_aeb_2_area:avs_rmap_0_read_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write                             : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write -> rmap_mem_ffee_aeb_2_area:avs_rmap_0_write_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata -> rmap_mem_ffee_aeb_2_area:avs_rmap_0_writedata_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata                          : std_logic_vector(31 downto 0);  -- rmap_mem_ffee_aeb_3_area:avs_rmap_0_readdata_o -> mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest                       : std_logic;                      -- rmap_mem_ffee_aeb_3_area:avs_rmap_0_waitrequest_o -> mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address -> rmap_mem_ffee_aeb_3_area:avs_rmap_0_address_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read                              : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read -> rmap_mem_ffee_aeb_3_area:avs_rmap_0_read_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write                             : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write -> rmap_mem_ffee_aeb_3_area:avs_rmap_0_write_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata -> rmap_mem_ffee_aeb_3_area:avs_rmap_0_writedata_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata                          : std_logic_vector(31 downto 0);  -- rmap_mem_ffee_aeb_4_area:avs_rmap_0_readdata_o -> mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest                       : std_logic;                      -- rmap_mem_ffee_aeb_4_area:avs_rmap_0_waitrequest_o -> mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address -> rmap_mem_ffee_aeb_4_area:avs_rmap_0_address_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read                              : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read -> rmap_mem_ffee_aeb_4_area:avs_rmap_0_read_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write                             : std_logic;                      -- mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write -> rmap_mem_ffee_aeb_4_area:avs_rmap_0_write_i
	signal mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata -> rmap_mem_ffee_aeb_4_area:avs_rmap_0_writedata_i
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_readdata                              : std_logic_vector(31 downto 0);  -- FTDI_UMFT601A_Module:avalon_slave_config_readdata_o -> mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_readdata
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_waitrequest                           : std_logic;                      -- FTDI_UMFT601A_Module:avalon_slave_config_waitrequest_o -> mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_waitrequest
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_address                               : std_logic_vector(7 downto 0);   -- mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_address -> FTDI_UMFT601A_Module:avalon_slave_config_address_i
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_read                                  : std_logic;                      -- mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_read -> FTDI_UMFT601A_Module:avalon_slave_config_read_i
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_write                                 : std_logic;                      -- mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_write -> FTDI_UMFT601A_Module:avalon_slave_config_write_i
	signal mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_writedata                             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:FTDI_UMFT601A_Module_avalon_slave_config_writedata -> FTDI_UMFT601A_Module:avalon_slave_config_writedata_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_readdata                                     : std_logic_vector(31 downto 0);  -- Memory_Filler:avalon_slave_config_readdata_o -> mm_interconnect_1:Memory_Filler_avalon_slave_config_readdata
	signal mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest                                  : std_logic;                      -- Memory_Filler:avalon_slave_config_waitrequest_o -> mm_interconnect_1:Memory_Filler_avalon_slave_config_waitrequest
	signal mm_interconnect_1_memory_filler_avalon_slave_config_address                                      : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Memory_Filler_avalon_slave_config_address -> Memory_Filler:avalon_slave_config_address_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_read                                         : std_logic;                      -- mm_interconnect_1:Memory_Filler_avalon_slave_config_read -> Memory_Filler:avalon_slave_config_read_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_byteenable                                   : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Memory_Filler_avalon_slave_config_byteenable -> Memory_Filler:avalon_slave_config_byteenable_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_write                                        : std_logic;                      -- mm_interconnect_1:Memory_Filler_avalon_slave_config_write -> Memory_Filler:avalon_slave_config_write_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_writedata                                    : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Memory_Filler_avalon_slave_config_writedata -> Memory_Filler:avalon_slave_config_writedata_i
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_readdata                                       : std_logic_vector(63 downto 0);  -- ddr2_address_span_extender:avs_cntl_readdata -> mm_interconnect_1:ddr2_address_span_extender_cntl_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_read                                           : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_read -> ddr2_address_span_extender:avs_cntl_read
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable                                     : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_cntl_byteenable -> ddr2_address_span_extender:avs_cntl_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_write                                          : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_write -> ddr2_address_span_extender:avs_cntl_write
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_writedata                                      : std_logic_vector(63 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_cntl_writedata -> ddr2_address_span_extender:avs_cntl_writedata
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata                                              : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address                                               : std_logic_vector(0 downto 0);   -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata                                          : std_logic_vector(31 downto 0);  -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest                                       : std_logic;                      -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess                                       : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address                                           : std_logic_vector(8 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read                                              : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable                                        : std_logic_vector(3 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write                                             : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdata                                                : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:s0_readdata -> mm_interconnect_1:clock_bridge_afi_50_s0_readdata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest                                             : std_logic;                      -- clock_bridge_afi_50:s0_waitrequest -> mm_interconnect_1:clock_bridge_afi_50_s0_waitrequest
	signal mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess                                             : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_debugaccess -> clock_bridge_afi_50:s0_debugaccess
	signal mm_interconnect_1_clock_bridge_afi_50_s0_address                                                 : std_logic_vector(11 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_address -> clock_bridge_afi_50:s0_address
	signal mm_interconnect_1_clock_bridge_afi_50_s0_read                                                    : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_read -> clock_bridge_afi_50:s0_read
	signal mm_interconnect_1_clock_bridge_afi_50_s0_byteenable                                              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_byteenable -> clock_bridge_afi_50:s0_byteenable
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid                                           : std_logic;                      -- clock_bridge_afi_50:s0_readdatavalid -> mm_interconnect_1:clock_bridge_afi_50_s0_readdatavalid
	signal mm_interconnect_1_clock_bridge_afi_50_s0_write                                                   : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_write -> clock_bridge_afi_50:s0_write
	signal mm_interconnect_1_clock_bridge_afi_50_s0_writedata                                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_writedata -> clock_bridge_afi_50:s0_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_burstcount                                              : std_logic_vector(0 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_burstcount -> clock_bridge_afi_50:s0_burstcount
	signal mm_interconnect_1_onchip_memory_s1_chipselect                                                    : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_1_onchip_memory_s1_readdata                                                      : std_logic_vector(31 downto 0);  -- onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	signal mm_interconnect_1_onchip_memory_s1_address                                                       : std_logic_vector(17 downto 0);  -- mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_1_onchip_memory_s1_byteenable                                                    : std_logic_vector(3 downto 0);   -- mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_1_onchip_memory_s1_write                                                         : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_1_onchip_memory_s1_writedata                                                     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_1_onchip_memory_s1_clken                                                         : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_1_ext_flash_uas_readdata                                                         : std_logic_vector(15 downto 0);  -- ext_flash:uas_readdata -> mm_interconnect_1:ext_flash_uas_readdata
	signal mm_interconnect_1_ext_flash_uas_waitrequest                                                      : std_logic;                      -- ext_flash:uas_waitrequest -> mm_interconnect_1:ext_flash_uas_waitrequest
	signal mm_interconnect_1_ext_flash_uas_debugaccess                                                      : std_logic;                      -- mm_interconnect_1:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	signal mm_interconnect_1_ext_flash_uas_address                                                          : std_logic_vector(25 downto 0);  -- mm_interconnect_1:ext_flash_uas_address -> ext_flash:uas_address
	signal mm_interconnect_1_ext_flash_uas_read                                                             : std_logic;                      -- mm_interconnect_1:ext_flash_uas_read -> ext_flash:uas_read
	signal mm_interconnect_1_ext_flash_uas_byteenable                                                       : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	signal mm_interconnect_1_ext_flash_uas_readdatavalid                                                    : std_logic;                      -- ext_flash:uas_readdatavalid -> mm_interconnect_1:ext_flash_uas_readdatavalid
	signal mm_interconnect_1_ext_flash_uas_lock                                                             : std_logic;                      -- mm_interconnect_1:ext_flash_uas_lock -> ext_flash:uas_lock
	signal mm_interconnect_1_ext_flash_uas_write                                                            : std_logic;                      -- mm_interconnect_1:ext_flash_uas_write -> ext_flash:uas_write
	signal mm_interconnect_1_ext_flash_uas_writedata                                                        : std_logic_vector(15 downto 0);  -- mm_interconnect_1:ext_flash_uas_writedata -> ext_flash:uas_writedata
	signal mm_interconnect_1_ext_flash_uas_burstcount                                                       : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata                             : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avs_s0_readdata -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest                          : std_logic;                      -- ddr2_address_span_extender:avs_s0_waitrequest -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_waitrequest
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address                              : std_logic_vector(28 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_address -> ddr2_address_span_extender:avs_s0_address
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read                                 : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_read -> ddr2_address_span_extender:avs_s0_read
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable                           : std_logic_vector(3 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_byteenable -> ddr2_address_span_extender:avs_s0_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid                        : std_logic;                      -- ddr2_address_span_extender:avs_s0_readdatavalid -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdatavalid
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write                                : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_write -> ddr2_address_span_extender:avs_s0_write
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_writedata -> ddr2_address_span_extender:avs_s0_writedata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount                           : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_burstcount -> ddr2_address_span_extender:avs_s0_burstcount
	signal clock_bridge_afi_50_m0_waitrequest                                                               : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_waitrequest -> clock_bridge_afi_50:m0_waitrequest
	signal clock_bridge_afi_50_m0_readdata                                                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_2:clock_bridge_afi_50_m0_readdata -> clock_bridge_afi_50:m0_readdata
	signal clock_bridge_afi_50_m0_debugaccess                                                               : std_logic;                      -- clock_bridge_afi_50:m0_debugaccess -> mm_interconnect_2:clock_bridge_afi_50_m0_debugaccess
	signal clock_bridge_afi_50_m0_address                                                                   : std_logic_vector(11 downto 0);  -- clock_bridge_afi_50:m0_address -> mm_interconnect_2:clock_bridge_afi_50_m0_address
	signal clock_bridge_afi_50_m0_read                                                                      : std_logic;                      -- clock_bridge_afi_50:m0_read -> mm_interconnect_2:clock_bridge_afi_50_m0_read
	signal clock_bridge_afi_50_m0_byteenable                                                                : std_logic_vector(3 downto 0);   -- clock_bridge_afi_50:m0_byteenable -> mm_interconnect_2:clock_bridge_afi_50_m0_byteenable
	signal clock_bridge_afi_50_m0_readdatavalid                                                             : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_readdatavalid -> clock_bridge_afi_50:m0_readdatavalid
	signal clock_bridge_afi_50_m0_writedata                                                                 : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:m0_writedata -> mm_interconnect_2:clock_bridge_afi_50_m0_writedata
	signal clock_bridge_afi_50_m0_write                                                                     : std_logic;                      -- clock_bridge_afi_50:m0_write -> mm_interconnect_2:clock_bridge_afi_50_m0_write
	signal clock_bridge_afi_50_m0_burstcount                                                                : std_logic_vector(0 downto 0);   -- clock_bridge_afi_50:m0_burstcount -> mm_interconnect_2:clock_bridge_afi_50_m0_burstcount
	signal mm_interconnect_2_sync_avalon_mm_slave_readdata                                                  : std_logic_vector(31 downto 0);  -- sync:avalon_slave_readdata_o -> mm_interconnect_2:sync_avalon_mm_slave_readdata
	signal mm_interconnect_2_sync_avalon_mm_slave_waitrequest                                               : std_logic;                      -- sync:avalon_slave_waitrequest_o -> mm_interconnect_2:sync_avalon_mm_slave_waitrequest
	signal mm_interconnect_2_sync_avalon_mm_slave_address                                                   : std_logic_vector(7 downto 0);   -- mm_interconnect_2:sync_avalon_mm_slave_address -> sync:avalon_slave_address_i
	signal mm_interconnect_2_sync_avalon_mm_slave_read                                                      : std_logic;                      -- mm_interconnect_2:sync_avalon_mm_slave_read -> sync:avalon_slave_read_i
	signal mm_interconnect_2_sync_avalon_mm_slave_write                                                     : std_logic;                      -- mm_interconnect_2:sync_avalon_mm_slave_write -> sync:avalon_slave_write_i
	signal mm_interconnect_2_sync_avalon_mm_slave_writedata                                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:sync_avalon_mm_slave_writedata -> sync:avalon_slave_writedata_i
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata                            : std_logic_vector(31 downto 0);  -- rst_controller:avalon_slave_rst_controller_readdata -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_readdata
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest                         : std_logic;                      -- rst_controller:avalon_slave_rst_controller_waitrequest -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_waitrequest
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address                             : std_logic_vector(3 downto 0);   -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_address -> rst_controller:avalon_slave_rst_controller_address
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read                                : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_read -> rst_controller:avalon_slave_rst_controller_read
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write                               : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_write -> rst_controller:avalon_slave_rst_controller_write
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata                           : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_writedata -> rst_controller:avalon_slave_rst_controller_writedata
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect            : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata              : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest           : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address               : std_logic_vector(7 downto 0);   -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read                  : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable            : std_logic_vector(3 downto 0);   -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write                 : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect                                                  : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_chipselect -> m1_ddr2_i2c_sda:chipselect
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata                                                    : std_logic_vector(31 downto 0);  -- m1_ddr2_i2c_sda:readdata -> mm_interconnect_2:m1_ddr2_i2c_sda_s1_readdata
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_address                                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_address -> m1_ddr2_i2c_sda:address
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_write                                                       : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_write -> mm_interconnect_2_m1_ddr2_i2c_sda_s1_write:in
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata                                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_writedata -> m1_ddr2_i2c_sda:writedata
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect                                                  : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_chipselect -> m1_ddr2_i2c_scl:chipselect
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata                                                    : std_logic_vector(31 downto 0);  -- m1_ddr2_i2c_scl:readdata -> mm_interconnect_2:m1_ddr2_i2c_scl_s1_readdata
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_address                                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_address -> m1_ddr2_i2c_scl:address
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_write                                                       : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_write -> mm_interconnect_2_m1_ddr2_i2c_scl_s1_write:in
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata                                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_writedata -> m1_ddr2_i2c_scl:writedata
	signal mm_interconnect_2_pio_button_s1_readdata                                                         : std_logic_vector(31 downto 0);  -- pio_BUTTON:readdata -> mm_interconnect_2:pio_BUTTON_s1_readdata
	signal mm_interconnect_2_pio_button_s1_address                                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_BUTTON_s1_address -> pio_BUTTON:address
	signal mm_interconnect_2_pio_led_s1_chipselect                                                          : std_logic;                      -- mm_interconnect_2:pio_LED_s1_chipselect -> pio_LED:chipselect
	signal mm_interconnect_2_pio_led_s1_readdata                                                            : std_logic_vector(31 downto 0);  -- pio_LED:readdata -> mm_interconnect_2:pio_LED_s1_readdata
	signal mm_interconnect_2_pio_led_s1_address                                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_LED_s1_address -> pio_LED:address
	signal mm_interconnect_2_pio_led_s1_write                                                               : std_logic;                      -- mm_interconnect_2:pio_LED_s1_write -> mm_interconnect_2_pio_led_s1_write:in
	signal mm_interconnect_2_pio_led_s1_writedata                                                           : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_LED_s1_writedata -> pio_LED:writedata
	signal mm_interconnect_2_timer_1ms_s1_chipselect                                                        : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_chipselect -> timer_1ms:chipselect
	signal mm_interconnect_2_timer_1ms_s1_readdata                                                          : std_logic_vector(15 downto 0);  -- timer_1ms:readdata -> mm_interconnect_2:timer_1ms_s1_readdata
	signal mm_interconnect_2_timer_1ms_s1_address                                                           : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1ms_s1_address -> timer_1ms:address
	signal mm_interconnect_2_timer_1ms_s1_write                                                             : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_write -> mm_interconnect_2_timer_1ms_s1_write:in
	signal mm_interconnect_2_timer_1ms_s1_writedata                                                         : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1ms_s1_writedata -> timer_1ms:writedata
	signal mm_interconnect_2_pio_dip_s1_readdata                                                            : std_logic_vector(31 downto 0);  -- pio_DIP:readdata -> mm_interconnect_2:pio_DIP_s1_readdata
	signal mm_interconnect_2_pio_dip_s1_address                                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_DIP_s1_address -> pio_DIP:address
	signal mm_interconnect_2_timer_1us_s1_chipselect                                                        : std_logic;                      -- mm_interconnect_2:timer_1us_s1_chipselect -> timer_1us:chipselect
	signal mm_interconnect_2_timer_1us_s1_readdata                                                          : std_logic_vector(15 downto 0);  -- timer_1us:readdata -> mm_interconnect_2:timer_1us_s1_readdata
	signal mm_interconnect_2_timer_1us_s1_address                                                           : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1us_s1_address -> timer_1us:address
	signal mm_interconnect_2_timer_1us_s1_write                                                             : std_logic;                      -- mm_interconnect_2:timer_1us_s1_write -> mm_interconnect_2_timer_1us_s1_write:in
	signal mm_interconnect_2_timer_1us_s1_writedata                                                         : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1us_s1_writedata -> timer_1us:writedata
	signal mm_interconnect_2_pio_ext_s1_readdata                                                            : std_logic_vector(31 downto 0);  -- pio_EXT:readdata -> mm_interconnect_2:pio_EXT_s1_readdata
	signal mm_interconnect_2_pio_ext_s1_address                                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_EXT_s1_address -> pio_EXT:address
	signal mm_interconnect_2_sd_card_wp_n_s1_readdata                                                       : std_logic_vector(31 downto 0);  -- sd_card_wp_n:readdata -> mm_interconnect_2:sd_card_wp_n_s1_readdata
	signal mm_interconnect_2_sd_card_wp_n_s1_address                                                        : std_logic_vector(1 downto 0);   -- mm_interconnect_2:sd_card_wp_n_s1_address -> sd_card_wp_n:address
	signal mm_interconnect_2_temp_scl_s1_chipselect                                                         : std_logic;                      -- mm_interconnect_2:temp_scl_s1_chipselect -> temp_scl:chipselect
	signal mm_interconnect_2_temp_scl_s1_readdata                                                           : std_logic_vector(31 downto 0);  -- temp_scl:readdata -> mm_interconnect_2:temp_scl_s1_readdata
	signal mm_interconnect_2_temp_scl_s1_address                                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_scl_s1_address -> temp_scl:address
	signal mm_interconnect_2_temp_scl_s1_write                                                              : std_logic;                      -- mm_interconnect_2:temp_scl_s1_write -> mm_interconnect_2_temp_scl_s1_write:in
	signal mm_interconnect_2_temp_scl_s1_writedata                                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_scl_s1_writedata -> temp_scl:writedata
	signal mm_interconnect_2_temp_sda_s1_chipselect                                                         : std_logic;                      -- mm_interconnect_2:temp_sda_s1_chipselect -> temp_sda:chipselect
	signal mm_interconnect_2_temp_sda_s1_readdata                                                           : std_logic_vector(31 downto 0);  -- temp_sda:readdata -> mm_interconnect_2:temp_sda_s1_readdata
	signal mm_interconnect_2_temp_sda_s1_address                                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_sda_s1_address -> temp_sda:address
	signal mm_interconnect_2_temp_sda_s1_write                                                              : std_logic;                      -- mm_interconnect_2:temp_sda_s1_write -> mm_interconnect_2_temp_sda_s1_write:in
	signal mm_interconnect_2_temp_sda_s1_writedata                                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_sda_s1_writedata -> temp_sda:writedata
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect                                                  : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_chipselect -> m2_ddr2_i2c_sda:chipselect
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata                                                    : std_logic_vector(31 downto 0);  -- m2_ddr2_i2c_sda:readdata -> mm_interconnect_2:m2_ddr2_i2c_sda_s1_readdata
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_address                                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_address -> m2_ddr2_i2c_sda:address
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_write                                                       : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_write -> mm_interconnect_2_m2_ddr2_i2c_sda_s1_write:in
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata                                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_writedata -> m2_ddr2_i2c_sda:writedata
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect                                                  : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_chipselect -> m2_ddr2_i2c_scl:chipselect
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata                                                    : std_logic_vector(31 downto 0);  -- m2_ddr2_i2c_scl:readdata -> mm_interconnect_2:m2_ddr2_i2c_scl_s1_readdata
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_address                                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_address -> m2_ddr2_i2c_scl:address
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_write                                                       : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_write -> mm_interconnect_2_m2_ddr2_i2c_scl_s1_write:in
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata                                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_writedata -> m2_ddr2_i2c_scl:writedata
	signal mm_interconnect_2_csense_sdo_s1_readdata                                                         : std_logic_vector(31 downto 0);  -- csense_sdo:readdata -> mm_interconnect_2:csense_sdo_s1_readdata
	signal mm_interconnect_2_csense_sdo_s1_address                                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdo_s1_address -> csense_sdo:address
	signal mm_interconnect_2_csense_sdi_s1_chipselect                                                       : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_chipselect -> csense_sdi:chipselect
	signal mm_interconnect_2_csense_sdi_s1_readdata                                                         : std_logic_vector(31 downto 0);  -- csense_sdi:readdata -> mm_interconnect_2:csense_sdi_s1_readdata
	signal mm_interconnect_2_csense_sdi_s1_address                                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdi_s1_address -> csense_sdi:address
	signal mm_interconnect_2_csense_sdi_s1_write                                                            : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_write -> mm_interconnect_2_csense_sdi_s1_write:in
	signal mm_interconnect_2_csense_sdi_s1_writedata                                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sdi_s1_writedata -> csense_sdi:writedata
	signal mm_interconnect_2_csense_sck_s1_chipselect                                                       : std_logic;                      -- mm_interconnect_2:csense_sck_s1_chipselect -> csense_sck:chipselect
	signal mm_interconnect_2_csense_sck_s1_readdata                                                         : std_logic_vector(31 downto 0);  -- csense_sck:readdata -> mm_interconnect_2:csense_sck_s1_readdata
	signal mm_interconnect_2_csense_sck_s1_address                                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sck_s1_address -> csense_sck:address
	signal mm_interconnect_2_csense_sck_s1_write                                                            : std_logic;                      -- mm_interconnect_2:csense_sck_s1_write -> mm_interconnect_2_csense_sck_s1_write:in
	signal mm_interconnect_2_csense_sck_s1_writedata                                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sck_s1_writedata -> csense_sck:writedata
	signal mm_interconnect_2_csense_cs_n_s1_chipselect                                                      : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_chipselect -> csense_cs_n:chipselect
	signal mm_interconnect_2_csense_cs_n_s1_readdata                                                        : std_logic_vector(31 downto 0);  -- csense_cs_n:readdata -> mm_interconnect_2:csense_cs_n_s1_readdata
	signal mm_interconnect_2_csense_cs_n_s1_address                                                         : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_cs_n_s1_address -> csense_cs_n:address
	signal mm_interconnect_2_csense_cs_n_s1_write                                                           : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_write -> mm_interconnect_2_csense_cs_n_s1_write:in
	signal mm_interconnect_2_csense_cs_n_s1_writedata                                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_cs_n_s1_writedata -> csense_cs_n:writedata
	signal mm_interconnect_2_csense_adc_fo_s1_chipselect                                                    : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_chipselect -> csense_adc_fo:chipselect
	signal mm_interconnect_2_csense_adc_fo_s1_readdata                                                      : std_logic_vector(31 downto 0);  -- csense_adc_fo:readdata -> mm_interconnect_2:csense_adc_fo_s1_readdata
	signal mm_interconnect_2_csense_adc_fo_s1_address                                                       : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_adc_fo_s1_address -> csense_adc_fo:address
	signal mm_interconnect_2_csense_adc_fo_s1_write                                                         : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_write -> mm_interconnect_2_csense_adc_fo_s1_write:in
	signal mm_interconnect_2_csense_adc_fo_s1_writedata                                                     : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_adc_fo_s1_writedata -> csense_adc_fo:writedata
	signal mm_interconnect_2_pio_led_painel_s1_chipselect                                                   : std_logic;                      -- mm_interconnect_2:pio_LED_painel_s1_chipselect -> pio_LED_painel:chipselect
	signal mm_interconnect_2_pio_led_painel_s1_readdata                                                     : std_logic_vector(31 downto 0);  -- pio_LED_painel:readdata -> mm_interconnect_2:pio_LED_painel_s1_readdata
	signal mm_interconnect_2_pio_led_painel_s1_address                                                      : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_LED_painel_s1_address -> pio_LED_painel:address
	signal mm_interconnect_2_pio_led_painel_s1_write                                                        : std_logic;                      -- mm_interconnect_2:pio_LED_painel_s1_write -> mm_interconnect_2_pio_led_painel_s1_write:in
	signal mm_interconnect_2_pio_led_painel_s1_writedata                                                    : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_LED_painel_s1_writedata -> pio_LED_painel:writedata
	signal mm_interconnect_2_rtcc_alarm_s1_readdata                                                         : std_logic_vector(31 downto 0);  -- rtcc_alarm:readdata -> mm_interconnect_2:rtcc_alarm_s1_readdata
	signal mm_interconnect_2_rtcc_alarm_s1_address                                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_alarm_s1_address -> rtcc_alarm:address
	signal mm_interconnect_2_rtcc_sdo_s1_readdata                                                           : std_logic_vector(31 downto 0);  -- rtcc_sdo:readdata -> mm_interconnect_2:rtcc_sdo_s1_readdata
	signal mm_interconnect_2_rtcc_sdo_s1_address                                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sdo_s1_address -> rtcc_sdo:address
	signal mm_interconnect_2_rtcc_sdi_s1_chipselect                                                         : std_logic;                      -- mm_interconnect_2:rtcc_sdi_s1_chipselect -> rtcc_sdi:chipselect
	signal mm_interconnect_2_rtcc_sdi_s1_readdata                                                           : std_logic_vector(31 downto 0);  -- rtcc_sdi:readdata -> mm_interconnect_2:rtcc_sdi_s1_readdata
	signal mm_interconnect_2_rtcc_sdi_s1_address                                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sdi_s1_address -> rtcc_sdi:address
	signal mm_interconnect_2_rtcc_sdi_s1_write                                                              : std_logic;                      -- mm_interconnect_2:rtcc_sdi_s1_write -> mm_interconnect_2_rtcc_sdi_s1_write:in
	signal mm_interconnect_2_rtcc_sdi_s1_writedata                                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_sdi_s1_writedata -> rtcc_sdi:writedata
	signal mm_interconnect_2_rtcc_sck_s1_chipselect                                                         : std_logic;                      -- mm_interconnect_2:rtcc_sck_s1_chipselect -> rtcc_sck:chipselect
	signal mm_interconnect_2_rtcc_sck_s1_readdata                                                           : std_logic_vector(31 downto 0);  -- rtcc_sck:readdata -> mm_interconnect_2:rtcc_sck_s1_readdata
	signal mm_interconnect_2_rtcc_sck_s1_address                                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sck_s1_address -> rtcc_sck:address
	signal mm_interconnect_2_rtcc_sck_s1_write                                                              : std_logic;                      -- mm_interconnect_2:rtcc_sck_s1_write -> mm_interconnect_2_rtcc_sck_s1_write:in
	signal mm_interconnect_2_rtcc_sck_s1_writedata                                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_sck_s1_writedata -> rtcc_sck:writedata
	signal mm_interconnect_2_rtcc_cs_n_s1_chipselect                                                        : std_logic;                      -- mm_interconnect_2:rtcc_cs_n_s1_chipselect -> rtcc_cs_n:chipselect
	signal mm_interconnect_2_rtcc_cs_n_s1_readdata                                                          : std_logic_vector(31 downto 0);  -- rtcc_cs_n:readdata -> mm_interconnect_2:rtcc_cs_n_s1_readdata
	signal mm_interconnect_2_rtcc_cs_n_s1_address                                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_cs_n_s1_address -> rtcc_cs_n:address
	signal mm_interconnect_2_rtcc_cs_n_s1_write                                                             : std_logic;                      -- mm_interconnect_2:rtcc_cs_n_s1_write -> mm_interconnect_2_rtcc_cs_n_s1_write:in
	signal mm_interconnect_2_rtcc_cs_n_s1_writedata                                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_cs_n_s1_writedata -> rtcc_cs_n:writedata
	signal mm_interconnect_2_rs232_uart_s1_chipselect                                                       : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_chipselect -> rs232_uart:chipselect
	signal mm_interconnect_2_rs232_uart_s1_readdata                                                         : std_logic_vector(15 downto 0);  -- rs232_uart:readdata -> mm_interconnect_2:rs232_uart_s1_readdata
	signal mm_interconnect_2_rs232_uart_s1_address                                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_2:rs232_uart_s1_address -> rs232_uart:address
	signal mm_interconnect_2_rs232_uart_s1_read                                                             : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_read -> mm_interconnect_2_rs232_uart_s1_read:in
	signal mm_interconnect_2_rs232_uart_s1_begintransfer                                                    : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_begintransfer -> rs232_uart:begintransfer
	signal mm_interconnect_2_rs232_uart_s1_write                                                            : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_write -> mm_interconnect_2_rs232_uart_s1_write:in
	signal mm_interconnect_2_rs232_uart_s1_writedata                                                        : std_logic_vector(15 downto 0);  -- mm_interconnect_2:rs232_uart_s1_writedata -> rs232_uart:writedata
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect                                                 : std_logic;                      -- mm_interconnect_2:pio_ctrl_io_lvds_s1_chipselect -> pio_ctrl_io_lvds:chipselect
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata                                                   : std_logic_vector(31 downto 0);  -- pio_ctrl_io_lvds:readdata -> mm_interconnect_2:pio_ctrl_io_lvds_s1_readdata
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_address                                                    : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_ctrl_io_lvds_s1_address -> pio_ctrl_io_lvds:address
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_write                                                      : std_logic;                      -- mm_interconnect_2:pio_ctrl_io_lvds_s1_write -> mm_interconnect_2_pio_ctrl_io_lvds_s1_write:in
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata                                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_ctrl_io_lvds_s1_writedata -> pio_ctrl_io_lvds:writedata
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_1_select_s1_chipselect -> pio_spw_demux_ch_1_select:chipselect
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_readdata                                          : std_logic_vector(31 downto 0);  -- pio_spw_demux_ch_1_select:readdata -> mm_interconnect_2:pio_spw_demux_ch_1_select_s1_readdata
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_spw_demux_ch_1_select_s1_address -> pio_spw_demux_ch_1_select:address
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write                                             : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_1_select_s1_write -> mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write:in
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_spw_demux_ch_1_select_s1_writedata -> pio_spw_demux_ch_1_select:writedata
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_2_select_s1_chipselect -> pio_spw_demux_ch_2_select:chipselect
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_readdata                                          : std_logic_vector(31 downto 0);  -- pio_spw_demux_ch_2_select:readdata -> mm_interconnect_2:pio_spw_demux_ch_2_select_s1_readdata
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_spw_demux_ch_2_select_s1_address -> pio_spw_demux_ch_2_select:address
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write                                             : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_2_select_s1_write -> mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write:in
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_spw_demux_ch_2_select_s1_writedata -> pio_spw_demux_ch_2_select:writedata
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_3_select_s1_chipselect -> pio_spw_demux_ch_3_select:chipselect
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_readdata                                          : std_logic_vector(31 downto 0);  -- pio_spw_demux_ch_3_select:readdata -> mm_interconnect_2:pio_spw_demux_ch_3_select_s1_readdata
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_spw_demux_ch_3_select_s1_address -> pio_spw_demux_ch_3_select:address
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write                                             : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_3_select_s1_write -> mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write:in
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_spw_demux_ch_3_select_s1_writedata -> pio_spw_demux_ch_3_select:writedata
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_4_select_s1_chipselect -> pio_spw_demux_ch_4_select:chipselect
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_readdata                                          : std_logic_vector(31 downto 0);  -- pio_spw_demux_ch_4_select:readdata -> mm_interconnect_2:pio_spw_demux_ch_4_select_s1_readdata
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_spw_demux_ch_4_select_s1_address -> pio_spw_demux_ch_4_select:address
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write                                             : std_logic;                      -- mm_interconnect_2:pio_spw_demux_ch_4_select_s1_write -> mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write:in
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_spw_demux_ch_4_select_s1_writedata -> pio_spw_demux_ch_4_select:writedata
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_chipselect                                   : std_logic;                      -- mm_interconnect_2:pio_ftdi_umft601a_module_reset_s1_chipselect -> pio_ftdi_umft601a_module_reset:chipselect
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_readdata                                     : std_logic_vector(31 downto 0);  -- pio_ftdi_umft601a_module_reset:readdata -> mm_interconnect_2:pio_ftdi_umft601a_module_reset_s1_readdata
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_address                                      : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_ftdi_umft601a_module_reset_s1_address -> pio_ftdi_umft601a_module_reset:address
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write                                        : std_logic;                      -- mm_interconnect_2:pio_ftdi_umft601a_module_reset_s1_write -> mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write:in
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_writedata                                    : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_ftdi_umft601a_module_reset_s1_writedata -> pio_ftdi_umft601a_module_reset:writedata
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_chipselect                                      : std_logic;                      -- mm_interconnect_2:pio_iso_logic_signal_enable_s1_chipselect -> pio_iso_logic_signal_enable:chipselect
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_readdata                                        : std_logic_vector(31 downto 0);  -- pio_iso_logic_signal_enable:readdata -> mm_interconnect_2:pio_iso_logic_signal_enable_s1_readdata
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_address                                         : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_iso_logic_signal_enable_s1_address -> pio_iso_logic_signal_enable:address
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_write                                           : std_logic;                      -- mm_interconnect_2:pio_iso_logic_signal_enable_s1_write -> mm_interconnect_2_pio_iso_logic_signal_enable_s1_write:in
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_iso_logic_signal_enable_s1_writedata -> pio_iso_logic_signal_enable:writedata
	signal m1_clock_bridge_m0_waitrequest                                                                   : std_logic;                      -- mm_interconnect_3:m1_clock_bridge_m0_waitrequest -> m1_clock_bridge:m0_waitrequest
	signal m1_clock_bridge_m0_readdata                                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_3:m1_clock_bridge_m0_readdata -> m1_clock_bridge:m0_readdata
	signal m1_clock_bridge_m0_debugaccess                                                                   : std_logic;                      -- m1_clock_bridge:m0_debugaccess -> mm_interconnect_3:m1_clock_bridge_m0_debugaccess
	signal m1_clock_bridge_m0_address                                                                       : std_logic_vector(30 downto 0);  -- m1_clock_bridge:m0_address -> mm_interconnect_3:m1_clock_bridge_m0_address
	signal m1_clock_bridge_m0_read                                                                          : std_logic;                      -- m1_clock_bridge:m0_read -> mm_interconnect_3:m1_clock_bridge_m0_read
	signal m1_clock_bridge_m0_byteenable                                                                    : std_logic_vector(31 downto 0);  -- m1_clock_bridge:m0_byteenable -> mm_interconnect_3:m1_clock_bridge_m0_byteenable
	signal m1_clock_bridge_m0_readdatavalid                                                                 : std_logic;                      -- mm_interconnect_3:m1_clock_bridge_m0_readdatavalid -> m1_clock_bridge:m0_readdatavalid
	signal m1_clock_bridge_m0_writedata                                                                     : std_logic_vector(255 downto 0); -- m1_clock_bridge:m0_writedata -> mm_interconnect_3:m1_clock_bridge_m0_writedata
	signal m1_clock_bridge_m0_write                                                                         : std_logic;                      -- m1_clock_bridge:m0_write -> mm_interconnect_3:m1_clock_bridge_m0_write
	signal m1_clock_bridge_m0_burstcount                                                                    : std_logic_vector(2 downto 0);   -- m1_clock_bridge:m0_burstcount -> mm_interconnect_3:m1_clock_bridge_m0_burstcount
	signal mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer                                          : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_beginbursttransfer -> m1_ddr2_memory:avl_burstbegin
	signal mm_interconnect_3_m1_ddr2_memory_avl_readdata                                                    : std_logic_vector(255 downto 0); -- m1_ddr2_memory:avl_rdata -> mm_interconnect_3:m1_ddr2_memory_avl_readdata
	signal m1_ddr2_memory_avl_waitrequest                                                                   : std_logic;                      -- m1_ddr2_memory:avl_ready -> m1_ddr2_memory_avl_waitrequest:in
	signal mm_interconnect_3_m1_ddr2_memory_avl_address                                                     : std_logic_vector(25 downto 0);  -- mm_interconnect_3:m1_ddr2_memory_avl_address -> m1_ddr2_memory:avl_addr
	signal mm_interconnect_3_m1_ddr2_memory_avl_read                                                        : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_read -> m1_ddr2_memory:avl_read_req
	signal mm_interconnect_3_m1_ddr2_memory_avl_byteenable                                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_3:m1_ddr2_memory_avl_byteenable -> m1_ddr2_memory:avl_be
	signal mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid                                               : std_logic;                      -- m1_ddr2_memory:avl_rdata_valid -> mm_interconnect_3:m1_ddr2_memory_avl_readdatavalid
	signal mm_interconnect_3_m1_ddr2_memory_avl_write                                                       : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_write -> m1_ddr2_memory:avl_write_req
	signal mm_interconnect_3_m1_ddr2_memory_avl_writedata                                                   : std_logic_vector(255 downto 0); -- mm_interconnect_3:m1_ddr2_memory_avl_writedata -> m1_ddr2_memory:avl_wdata
	signal mm_interconnect_3_m1_ddr2_memory_avl_burstcount                                                  : std_logic_vector(7 downto 0);   -- mm_interconnect_3:m1_ddr2_memory_avl_burstcount -> m1_ddr2_memory:avl_size
	signal m1_ddr2_memory_afi_clk_clk                                                                       : std_logic;                      -- m1_ddr2_memory:afi_clk -> [mm_interconnect_3:m1_ddr2_memory_afi_clk_clk, rst_controller_008:clk]
	signal irq_mapper_receiver0_irq                                                                         : std_logic;                      -- Communication_Module_v2_Ch1:feeb_interrupt_sender_irq_o -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                         : std_logic;                      -- Communication_Module_v2_Ch2:feeb_interrupt_sender_irq_o -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                         : std_logic;                      -- Communication_Module_v2_Ch4:feeb_interrupt_sender_irq_o -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                         : std_logic;                      -- Communication_Module_v2_Ch3:feeb_interrupt_sender_irq_o -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                         : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver9_irq                                                                         : std_logic;                      -- Communication_Module_v2_Ch1:rmap_interrupt_sender_irq_o -> irq_mapper:receiver9_irq
	signal irq_mapper_receiver10_irq                                                                        : std_logic;                      -- Communication_Module_v2_Ch2:rmap_interrupt_sender_irq_o -> irq_mapper:receiver10_irq
	signal irq_mapper_receiver11_irq                                                                        : std_logic;                      -- Communication_Module_v2_Ch4:rmap_interrupt_sender_irq_o -> irq_mapper:receiver11_irq
	signal irq_mapper_receiver12_irq                                                                        : std_logic;                      -- Communication_Module_v2_Ch3:rmap_interrupt_sender_irq_o -> irq_mapper:receiver12_irq
	signal irq_mapper_receiver13_irq                                                                        : std_logic;                      -- FTDI_UMFT601A_Module:rx_interrupt_sender_irq_o -> irq_mapper:receiver13_irq
	signal irq_mapper_receiver15_irq                                                                        : std_logic;                      -- FTDI_UMFT601A_Module:tx_interrupt_sender_irq_o -> irq_mapper:receiver15_irq
	signal nios2_gen2_0_irq_irq                                                                             : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver5_irq                                                                         : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver5_irq
	signal irq_synchronizer_receiver_irq                                                                    : std_logic_vector(0 downto 0);   -- timer_1ms:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver6_irq                                                                         : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver6_irq
	signal irq_synchronizer_001_receiver_irq                                                                : std_logic_vector(0 downto 0);   -- timer_1us:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver7_irq                                                                         : std_logic;                      -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver7_irq
	signal irq_synchronizer_002_receiver_irq                                                                : std_logic_vector(0 downto 0);   -- rs232_uart:irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver8_irq                                                                         : std_logic;                      -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver8_irq
	signal irq_synchronizer_003_receiver_irq                                                                : std_logic_vector(0 downto 0);   -- sync:pre_sync_interrupt_sender_irq_o -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver14_irq                                                                        : std_logic;                      -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver14_irq
	signal irq_synchronizer_004_receiver_irq                                                                : std_logic_vector(0 downto 0);   -- sync:sync_interrupt_sender_irq_o -> irq_synchronizer_004:receiver_irq
	signal rst_controller_001_reset_out_reset                                                               : std_logic;                      -- rst_controller_001:reset_out -> [clock_bridge_afi_50:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, mm_interconnect_2:clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset, rst_controller:reset_sink_reset, rst_controller_001_reset_out_reset:in, sync:reset_sink_reset_i]
	signal rst_controller_002_reset_out_reset                                                               : std_logic;                      -- rst_controller_002:reset_out -> [Communication_Module_v2_Ch1:reset_sink_reset_i, Communication_Module_v2_Ch2:reset_sink_reset_i, Communication_Module_v2_Ch3:reset_sink_reset_i, Communication_Module_v2_Ch4:reset_sink_reset_i, FTDI_UMFT601A_Module:reset_sink_reset_i, Memory_Filler:reset_sink_reset_i, SpaceWire_Demux_Ch1:reset_i, SpaceWire_Demux_Ch2:reset_i, SpaceWire_Demux_Ch3:reset_i, SpaceWire_Demux_Ch4:reset_i, clock_bridge_afi_50:s0_reset, ddr2_address_span_extender:reset, m1_clock_bridge:s0_reset, mm_interconnect_0:FTDI_UMFT601A_Module_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rmap_mem_ffee_aeb_1_area:reset_i, rmap_mem_ffee_aeb_2_area:reset_i, rmap_mem_ffee_aeb_3_area:reset_i, rmap_mem_ffee_aeb_4_area:reset_i, rmap_mem_ffee_deb_area:reset_i, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                                                           : std_logic;                      -- rst_controller_002:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	signal rst_controller_003_reset_out_reset                                                               : std_logic;                      -- rst_controller_003:reset_out -> [SpaceWire_Channel_A:reset_i, SpaceWire_Channel_B:reset_i, SpaceWire_Channel_C:reset_i, SpaceWire_Channel_D:reset_i, SpaceWire_Channel_E:reset_i, SpaceWire_Channel_F:reset_i, SpaceWire_Channel_G:reset_i, SpaceWire_Channel_H:reset_i, mm_interconnect_0:m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]
	signal rst_controller_004_reset_out_reset                                                               : std_logic;                      -- rst_controller_004:reset_out -> [ext_flash:reset_reset, mm_interconnect_1:ext_flash_reset_reset_bridge_in_reset_reset, tristate_conduit_bridge_0:reset]
	signal rst_controller_005_reset_out_reset                                                               : std_logic;                      -- rst_controller_005:reset_out -> [m1_clock_bridge:m0_reset, mm_interconnect_3:m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_006_reset_out_reset                                                               : std_logic;                      -- rst_controller_006:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_006_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_006_reset_out_reset_req                                                           : std_logic;                      -- rst_controller_006:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_007_reset_out_reset                                                               : std_logic;                      -- rst_controller_007:reset_out -> [irq_synchronizer_002:receiver_reset, mm_interconnect_2:rs232_uart_reset_reset_bridge_in_reset_reset, rst_controller_007_reset_out_reset:in]
	signal rst_controller_reset_source_rs232_reset                                                          : std_logic;                      -- rst_controller:reset_source_rs232_reset -> rst_controller_007:reset_in1
	signal rst_controller_008_reset_out_reset                                                               : std_logic;                      -- rst_controller_008:reset_out -> [mm_interconnect_3:m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]
	signal rst_reset_n_ports_inv                                                                            : std_logic;                      -- rst_reset_n:inv -> [rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_004:reset_in1, rst_controller_005:reset_in0, rst_controller_006:reset_in0, rst_controller_007:reset_in0, rst_controller_008:reset_in0]
	signal mm_interconnect_0_m2_ddr2_memory_avl_inv                                                         : std_logic;                      -- m2_ddr2_memory_avl_waitrequest:inv -> mm_interconnect_0:m2_ddr2_memory_avl_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv                                   : std_logic;                      -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv                                  : std_logic;                      -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv                                             : std_logic;                      -- mm_interconnect_2_m1_ddr2_i2c_sda_s1_write:inv -> m1_ddr2_i2c_sda:write_n
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv                                             : std_logic;                      -- mm_interconnect_2_m1_ddr2_i2c_scl_s1_write:inv -> m1_ddr2_i2c_scl:write_n
	signal mm_interconnect_2_pio_led_s1_write_ports_inv                                                     : std_logic;                      -- mm_interconnect_2_pio_led_s1_write:inv -> pio_LED:write_n
	signal mm_interconnect_2_timer_1ms_s1_write_ports_inv                                                   : std_logic;                      -- mm_interconnect_2_timer_1ms_s1_write:inv -> timer_1ms:write_n
	signal mm_interconnect_2_timer_1us_s1_write_ports_inv                                                   : std_logic;                      -- mm_interconnect_2_timer_1us_s1_write:inv -> timer_1us:write_n
	signal mm_interconnect_2_temp_scl_s1_write_ports_inv                                                    : std_logic;                      -- mm_interconnect_2_temp_scl_s1_write:inv -> temp_scl:write_n
	signal mm_interconnect_2_temp_sda_s1_write_ports_inv                                                    : std_logic;                      -- mm_interconnect_2_temp_sda_s1_write:inv -> temp_sda:write_n
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv                                             : std_logic;                      -- mm_interconnect_2_m2_ddr2_i2c_sda_s1_write:inv -> m2_ddr2_i2c_sda:write_n
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv                                             : std_logic;                      -- mm_interconnect_2_m2_ddr2_i2c_scl_s1_write:inv -> m2_ddr2_i2c_scl:write_n
	signal mm_interconnect_2_csense_sdi_s1_write_ports_inv                                                  : std_logic;                      -- mm_interconnect_2_csense_sdi_s1_write:inv -> csense_sdi:write_n
	signal mm_interconnect_2_csense_sck_s1_write_ports_inv                                                  : std_logic;                      -- mm_interconnect_2_csense_sck_s1_write:inv -> csense_sck:write_n
	signal mm_interconnect_2_csense_cs_n_s1_write_ports_inv                                                 : std_logic;                      -- mm_interconnect_2_csense_cs_n_s1_write:inv -> csense_cs_n:write_n
	signal mm_interconnect_2_csense_adc_fo_s1_write_ports_inv                                               : std_logic;                      -- mm_interconnect_2_csense_adc_fo_s1_write:inv -> csense_adc_fo:write_n
	signal mm_interconnect_2_pio_led_painel_s1_write_ports_inv                                              : std_logic;                      -- mm_interconnect_2_pio_led_painel_s1_write:inv -> pio_LED_painel:write_n
	signal mm_interconnect_2_rtcc_sdi_s1_write_ports_inv                                                    : std_logic;                      -- mm_interconnect_2_rtcc_sdi_s1_write:inv -> rtcc_sdi:write_n
	signal mm_interconnect_2_rtcc_sck_s1_write_ports_inv                                                    : std_logic;                      -- mm_interconnect_2_rtcc_sck_s1_write:inv -> rtcc_sck:write_n
	signal mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv                                                   : std_logic;                      -- mm_interconnect_2_rtcc_cs_n_s1_write:inv -> rtcc_cs_n:write_n
	signal mm_interconnect_2_rs232_uart_s1_read_ports_inv                                                   : std_logic;                      -- mm_interconnect_2_rs232_uart_s1_read:inv -> rs232_uart:read_n
	signal mm_interconnect_2_rs232_uart_s1_write_ports_inv                                                  : std_logic;                      -- mm_interconnect_2_rs232_uart_s1_write:inv -> rs232_uart:write_n
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv                                            : std_logic;                      -- mm_interconnect_2_pio_ctrl_io_lvds_s1_write:inv -> pio_ctrl_io_lvds:write_n
	signal mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write:inv -> pio_spw_demux_ch_1_select:write_n
	signal mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write:inv -> pio_spw_demux_ch_2_select:write_n
	signal mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write:inv -> pio_spw_demux_ch_3_select:write_n
	signal mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write:inv -> pio_spw_demux_ch_4_select:write_n
	signal mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write_ports_inv                              : std_logic;                      -- mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write:inv -> pio_ftdi_umft601a_module_reset:write_n
	signal mm_interconnect_2_pio_iso_logic_signal_enable_s1_write_ports_inv                                 : std_logic;                      -- mm_interconnect_2_pio_iso_logic_signal_enable_s1_write:inv -> pio_iso_logic_signal_enable:write_n
	signal mm_interconnect_3_m1_ddr2_memory_avl_inv                                                         : std_logic;                      -- m1_ddr2_memory_avl_waitrequest:inv -> mm_interconnect_3:m1_ddr2_memory_avl_waitrequest
	signal rst_controller_001_reset_out_reset_ports_inv                                                     : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, csense_adc_fo:reset_n, csense_cs_n:reset_n, csense_sck:reset_n, csense_sdi:reset_n, csense_sdo:reset_n, m1_ddr2_i2c_scl:reset_n, m1_ddr2_i2c_sda:reset_n, m2_ddr2_i2c_scl:reset_n, m2_ddr2_i2c_sda:reset_n, pio_BUTTON:reset_n, pio_DIP:reset_n, pio_EXT:reset_n, pio_LED:reset_n, pio_LED_painel:reset_n, pio_ctrl_io_lvds:reset_n, pio_ftdi_umft601a_module_reset:reset_n, pio_iso_logic_signal_enable:reset_n, pio_spw_demux_ch_1_select:reset_n, pio_spw_demux_ch_2_select:reset_n, pio_spw_demux_ch_3_select:reset_n, pio_spw_demux_ch_4_select:reset_n, rtcc_alarm:reset_n, rtcc_cs_n:reset_n, rtcc_sck:reset_n, rtcc_sdi:reset_n, rtcc_sdo:reset_n, sd_card_wp_n:reset_n, temp_scl:reset_n, temp_sda:reset_n, timer_1ms:reset_n, timer_1us:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                                                     : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> [jtag_uart_0:rst_n, sysid_qsys:reset_n]
	signal rst_controller_006_reset_out_reset_ports_inv                                                     : std_logic;                      -- rst_controller_006_reset_out_reset:inv -> nios2_gen2_0:reset_n
	signal rst_controller_007_reset_out_reset_ports_inv                                                     : std_logic;                      -- rst_controller_007_reset_out_reset:inv -> rs232_uart:reset_n

begin

	altera_up_sd_card_avalon_interface_0 : component Altera_UP_SD_Card_Avalon_Interface
		port map (
			i_avalon_chip_select => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  -- avalon_sdcard_slave.chipselect
			i_avalon_address     => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     --                    .address
			i_avalon_read        => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                    .read
			i_avalon_write       => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                    .write
			i_avalon_byteenable  => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                    .byteenable
			i_avalon_writedata   => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                    .writedata
			o_avalon_readdata    => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                    .readdata
			o_avalon_waitrequest => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                    .waitrequest
			i_clock              => clk50_clk,                                                                              --                 clk.clk
			i_reset_n            => rst_controller_001_reset_out_reset_ports_inv,                                           --               reset.reset_n
			b_SD_cmd             => sd_card_ip_b_SD_cmd,                                                                    --         conduit_end.export
			b_SD_dat             => sd_card_ip_b_SD_dat,                                                                    --                    .export
			b_SD_dat3            => sd_card_ip_b_SD_dat3,                                                                   --                    .export
			o_SD_clock           => sd_card_ip_o_SD_clock                                                                   --                    .export
		);

	communication_module_v2_ch1 : component comm_v2_top
		port map (
			reset_sink_reset_i                     => rst_controller_002_reset_out_reset,                                                               --                                   reset_sink.reset
			clock_sink_clk_i                       => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                                   clock_sink.clk
			channel_sync_i                         => comm_1_sync_sync_signal,                                                                          --                     conduit_end_channel_sync.sync_signal
			avs_config_address_i                   => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_address,                     --                       avalon_mm_config_slave.address
			avs_config_write_i                     => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_write,                       --                                             .write
			avs_config_writedata_i                 => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_writedata,                   --                                             .writedata
			avs_config_read_i                      => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_read,                        --                                             .read
			avs_config_readdata_o                  => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_readdata,                    --                                             .readdata
			avs_config_waitrequest_o               => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_waitrequest,                 --                                             .waitrequest
			avm_left_buffer_readdata_i             => communication_module_v2_ch1_avalon_mm_left_buffer_master_readdata,                                --                 avalon_mm_left_buffer_master.readdata
			avm_left_buffer_waitrequest_i          => communication_module_v2_ch1_avalon_mm_left_buffer_master_waitrequest,                             --                                             .waitrequest
			avm_left_buffer_address_o              => communication_module_v2_ch1_avalon_mm_left_buffer_master_address,                                 --                                             .address
			avm_left_buffer_read_o                 => communication_module_v2_ch1_avalon_mm_left_buffer_master_read,                                    --                                             .read
			avm_right_buffer_readdata_i            => communication_module_v2_ch1_avalon_mm_right_buffer_master_readdata,                               --                avalon_mm_right_buffer_master.readdata
			avm_right_buffer_waitrequest_i         => communication_module_v2_ch1_avalon_mm_right_buffer_master_waitrequest,                            --                                             .waitrequest
			avm_right_buffer_address_o             => communication_module_v2_ch1_avalon_mm_right_buffer_master_address,                                --                                             .address
			avm_right_buffer_read_o                => communication_module_v2_ch1_avalon_mm_right_buffer_master_read,                                   --                                             .read
			feeb_interrupt_sender_irq_o            => irq_mapper_receiver0_irq,                                                                         --                        feeb_interrupt_sender.irq
			rmap_interrupt_sender_irq_o            => irq_mapper_receiver9_irq,                                                                         --                        rmap_interrupt_sender.irq
			spw_link_status_started_i              => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --             conduit_end_spacewire_controller.spw_link_status_started_signal
			spw_link_status_connecting_i           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                             .spw_link_status_connecting_signal
			spw_link_status_running_i              => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                             .spw_link_status_running_signal
			spw_link_error_errdisc_i               => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                             .spw_link_error_errdisc_signal
			spw_link_error_errpar_i                => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                             .spw_link_error_errpar_signal
			spw_link_error_erresc_i                => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                             .spw_link_error_erresc_signal
			spw_link_error_errcred_i               => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                             .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_i             => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                             .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_i             => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                             .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_i             => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                             .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_i           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                             .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_i           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                             .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_i            => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                             .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_i            => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                             .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_i             => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                             .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_i           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                             .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_i          => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                             .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_i         => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                             .spw_errinj_ctrl_errinj_ready_signal
			spw_link_command_enable_o              => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --                                             .spw_link_command_enable_signal
			spw_link_command_autostart_o           => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                             .spw_link_command_autostart_signal
			spw_link_command_linkstart_o           => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                             .spw_link_command_linkstart_signal
			spw_link_command_linkdis_o             => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                             .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_o            => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                             .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_o              => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                             .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_o              => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                             .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_o              => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                             .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_o           => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                             .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_o          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                             .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_o           => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                             .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_o           => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                             .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_o         => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                             .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_o         => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                             .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_o          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                             .spw_errinj_ctrl_errinj_code_signal
			rmap_echo_echo_en_o                    => communication_module_v2_ch1_conduit_end_rmap_echo_out_echo_en_signal,                             --                    conduit_end_rmap_echo_out.echo_en_signal
			rmap_echo_echo_id_en_o                 => communication_module_v2_ch1_conduit_end_rmap_echo_out_echo_id_en_signal,                          --                                             .echo_id_en_signal
			rmap_echo_in_fifo_wrflag_o             => communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                      --                                             .in_fifo_wrflag_signal
			rmap_echo_in_fifo_wrdata_o             => communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                      --                                             .in_fifo_wrdata_signal
			rmap_echo_in_fifo_wrreq_o              => communication_module_v2_ch1_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                       --                                             .in_fifo_wrreq_signal
			rmap_echo_out_fifo_wrflag_o            => communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                     --                                             .out_fifo_wrflag_signal
			rmap_echo_out_fifo_wrdata_o            => communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                     --                                             .out_fifo_wrdata_signal
			rmap_echo_out_fifo_wrreq_o             => communication_module_v2_ch1_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                      --                                             .out_fifo_wrreq_signal
			rmm_deb_rmap_target_wr_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                        --  conduit_end_rmap_mem_deb_master_rmap_target.wr_waitrequest_signal
			rmm_deb_rmap_target_readdata_i         => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_rmap_target_rd_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_rmap_target_wr_address_o       => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal,        --                                             .wr_address_signal
			rmm_deb_rmap_target_write_o            => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,             --                                             .write_signal
			rmm_deb_rmap_target_writedata_o        => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,         --                                             .writedata_signal
			rmm_deb_rmap_target_rd_address_o       => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal,        --                                             .rd_address_signal
			rmm_deb_rmap_target_read_o             => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,              --                                             .read_signal
			rmm_deb_fee_hk_wr_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                        --       conduit_end_rmap_mem_deb_master_fee_hk.wr_waitrequest_signal
			rmm_deb_fee_hk_readdata_i              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_fee_hk_rd_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_fee_hk_wr_address_o            => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,             --                                             .wr_address_signal
			rmm_deb_fee_hk_write_o                 => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,                  --                                             .write_signal
			rmm_deb_fee_hk_writedata_o             => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,              --                                             .writedata_signal
			rmm_deb_fee_hk_rd_address_o            => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,             --                                             .rd_address_signal
			rmm_deb_fee_hk_read_o                  => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,                   --                                             .read_signal
			rmm_aeb1_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb1_master_rmap_target.wr_waitrequest_signal
			rmm_aeb1_rmap_target_readdata_i        => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_rmap_target_wr_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb1_rmap_target_write_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb1_rmap_target_writedata_o       => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb1_rmap_target_rd_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb1_rmap_target_read_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb1_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb1_master_fee_hk.wr_waitrequest_signal
			rmm_aeb1_fee_hk_readdata_i             => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_fee_hk_wr_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb1_fee_hk_write_o                => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb1_fee_hk_writedata_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb1_fee_hk_rd_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb1_fee_hk_read_o                 => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb2_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb2_master_rmap_target.wr_waitrequest_signal
			rmm_aeb2_rmap_target_readdata_i        => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_rmap_target_wr_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb2_rmap_target_write_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb2_rmap_target_writedata_o       => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb2_rmap_target_rd_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb2_rmap_target_read_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb2_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb2_master_fee_hk.wr_waitrequest_signal
			rmm_aeb2_fee_hk_readdata_i             => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_fee_hk_wr_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb2_fee_hk_write_o                => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb2_fee_hk_writedata_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb2_fee_hk_rd_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb2_fee_hk_read_o                 => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb3_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb3_master_rmap_target.wr_waitrequest_signal
			rmm_aeb3_rmap_target_readdata_i        => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_rmap_target_wr_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb3_rmap_target_write_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb3_rmap_target_writedata_o       => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb3_rmap_target_rd_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb3_rmap_target_read_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb3_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb3_master_fee_hk.wr_waitrequest_signal
			rmm_aeb3_fee_hk_readdata_i             => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_fee_hk_wr_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb3_fee_hk_write_o                => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb3_fee_hk_writedata_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb3_fee_hk_rd_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb3_fee_hk_read_o                 => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb4_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb4_master_rmap_target.wr_waitrequest_signal
			rmm_aeb4_rmap_target_readdata_i        => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_rmap_target_wr_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb4_rmap_target_write_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb4_rmap_target_writedata_o       => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb4_rmap_target_rd_address_o      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb4_rmap_target_read_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb4_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb4_master_fee_hk.wr_waitrequest_signal
			rmm_aeb4_fee_hk_readdata_i             => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_fee_hk_wr_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb4_fee_hk_write_o                => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb4_fee_hk_writedata_o            => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb4_fee_hk_rd_address_o           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb4_fee_hk_read_o                 => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,                  --                                             .read_signal
			channel_hk_rmap_target_status_o        => communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_status_signal,                 --                   conduit_end_channel_hk_out.rmap_target_status_signal
			channel_hk_rmap_target_indicate_o      => communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_indicate_signal,               --                                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_escape_err_signal,                --                                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_credit_err_signal,                --                                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_parity_err_signal,                --                                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_disconnect_signal,                --                                             .spw_link_disconnect_signal
			channel_hk_spw_link_started_o          => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_started_signal,                   --                                             .spw_link_started_signal
			channel_hk_spw_link_connecting_o       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_connecting_signal,                --                                             .spw_link_connecting_signal
			channel_hk_spw_link_running_o          => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_running_signal,                   --                                             .spw_link_running_signal
			channel_hk_frame_counter_o             => communication_module_v2_ch1_conduit_end_channel_hk_out_frame_counter_signal,                      --                                             .frame_counter_signal
			channel_hk_left_buffer_ccd_number_o    => communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,             --                                             .left_buffer_ccd_number_signal
			channel_hk_right_buffer_ccd_number_o   => communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,            --                                             .right_buffer_ccd_number_signal
			channel_hk_left_buffer_ccd_side_o      => communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,               --                                             .left_buffer_ccd_side_signal
			channel_hk_right_buffer_ccd_side_o     => communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,              --                                             .right_buffer_ccd_side_signal
			channel_hk_err_left_buffer_overflow_o  => communication_module_v2_ch1_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,           --                                             .err_left_buffer_overflow_signal
			channel_hk_err_right_buffer_overflow_o => communication_module_v2_ch1_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,          --                                             .err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_o          => communication_module_v2_ch1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal,          --             conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
			comm_data_control_data_hold_i          => comm_1_data_control_data_hold_signal,                                                             --                            comm_data_control.data_hold_signal
			comm_measurements_o                    => comm_1_measurements_measurements_signal                                                           --                conduit_end_comm_measurements.measurements_signal
		);

	communication_module_v2_ch2 : component comm_v2_top
		port map (
			reset_sink_reset_i                     => rst_controller_002_reset_out_reset,                                                               --                                   reset_sink.reset
			clock_sink_clk_i                       => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                                   clock_sink.clk
			channel_sync_i                         => comm_2_sync_sync_signal,                                                                          --                     conduit_end_channel_sync.sync_signal
			avs_config_address_i                   => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_address,                     --                       avalon_mm_config_slave.address
			avs_config_write_i                     => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_write,                       --                                             .write
			avs_config_writedata_i                 => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_writedata,                   --                                             .writedata
			avs_config_read_i                      => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_read,                        --                                             .read
			avs_config_readdata_o                  => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_readdata,                    --                                             .readdata
			avs_config_waitrequest_o               => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_waitrequest,                 --                                             .waitrequest
			avm_left_buffer_readdata_i             => communication_module_v2_ch2_avalon_mm_left_buffer_master_readdata,                                --                 avalon_mm_left_buffer_master.readdata
			avm_left_buffer_waitrequest_i          => communication_module_v2_ch2_avalon_mm_left_buffer_master_waitrequest,                             --                                             .waitrequest
			avm_left_buffer_address_o              => communication_module_v2_ch2_avalon_mm_left_buffer_master_address,                                 --                                             .address
			avm_left_buffer_read_o                 => communication_module_v2_ch2_avalon_mm_left_buffer_master_read,                                    --                                             .read
			avm_right_buffer_readdata_i            => communication_module_v2_ch2_avalon_mm_right_buffer_master_readdata,                               --                avalon_mm_right_buffer_master.readdata
			avm_right_buffer_waitrequest_i         => communication_module_v2_ch2_avalon_mm_right_buffer_master_waitrequest,                            --                                             .waitrequest
			avm_right_buffer_address_o             => communication_module_v2_ch2_avalon_mm_right_buffer_master_address,                                --                                             .address
			avm_right_buffer_read_o                => communication_module_v2_ch2_avalon_mm_right_buffer_master_read,                                   --                                             .read
			feeb_interrupt_sender_irq_o            => irq_mapper_receiver1_irq,                                                                         --                        feeb_interrupt_sender.irq
			rmap_interrupt_sender_irq_o            => irq_mapper_receiver10_irq,                                                                        --                        rmap_interrupt_sender.irq
			spw_link_status_started_i              => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --             conduit_end_spacewire_controller.spw_link_status_started_signal
			spw_link_status_connecting_i           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                             .spw_link_status_connecting_signal
			spw_link_status_running_i              => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                             .spw_link_status_running_signal
			spw_link_error_errdisc_i               => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                             .spw_link_error_errdisc_signal
			spw_link_error_errpar_i                => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                             .spw_link_error_errpar_signal
			spw_link_error_erresc_i                => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                             .spw_link_error_erresc_signal
			spw_link_error_errcred_i               => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                             .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_i             => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                             .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_i             => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                             .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_i             => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                             .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_i           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                             .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_i           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                             .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_i            => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                             .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_i            => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                             .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_i             => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                             .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_i           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                             .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_i          => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                             .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_i         => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                             .spw_errinj_ctrl_errinj_ready_signal
			spw_link_command_enable_o              => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --                                             .spw_link_command_enable_signal
			spw_link_command_autostart_o           => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                             .spw_link_command_autostart_signal
			spw_link_command_linkstart_o           => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                             .spw_link_command_linkstart_signal
			spw_link_command_linkdis_o             => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                             .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_o            => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                             .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_o              => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                             .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_o              => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                             .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_o              => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                             .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_o           => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                             .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_o          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                             .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_o           => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                             .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_o           => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                             .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_o         => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                             .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_o         => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                             .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_o          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                             .spw_errinj_ctrl_errinj_code_signal
			rmap_echo_echo_en_o                    => communication_module_v2_ch2_conduit_end_rmap_echo_out_echo_en_signal,                             --                    conduit_end_rmap_echo_out.echo_en_signal
			rmap_echo_echo_id_en_o                 => communication_module_v2_ch2_conduit_end_rmap_echo_out_echo_id_en_signal,                          --                                             .echo_id_en_signal
			rmap_echo_in_fifo_wrflag_o             => communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                      --                                             .in_fifo_wrflag_signal
			rmap_echo_in_fifo_wrdata_o             => communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                      --                                             .in_fifo_wrdata_signal
			rmap_echo_in_fifo_wrreq_o              => communication_module_v2_ch2_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                       --                                             .in_fifo_wrreq_signal
			rmap_echo_out_fifo_wrflag_o            => communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                     --                                             .out_fifo_wrflag_signal
			rmap_echo_out_fifo_wrdata_o            => communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                     --                                             .out_fifo_wrdata_signal
			rmap_echo_out_fifo_wrreq_o             => communication_module_v2_ch2_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                      --                                             .out_fifo_wrreq_signal
			rmm_deb_rmap_target_wr_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                        --  conduit_end_rmap_mem_deb_master_rmap_target.wr_waitrequest_signal
			rmm_deb_rmap_target_readdata_i         => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_rmap_target_rd_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_rmap_target_wr_address_o       => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal,        --                                             .wr_address_signal
			rmm_deb_rmap_target_write_o            => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,             --                                             .write_signal
			rmm_deb_rmap_target_writedata_o        => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,         --                                             .writedata_signal
			rmm_deb_rmap_target_rd_address_o       => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal,        --                                             .rd_address_signal
			rmm_deb_rmap_target_read_o             => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,              --                                             .read_signal
			rmm_deb_fee_hk_wr_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                        --       conduit_end_rmap_mem_deb_master_fee_hk.wr_waitrequest_signal
			rmm_deb_fee_hk_readdata_i              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_fee_hk_rd_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_fee_hk_wr_address_o            => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,             --                                             .wr_address_signal
			rmm_deb_fee_hk_write_o                 => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,                  --                                             .write_signal
			rmm_deb_fee_hk_writedata_o             => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,              --                                             .writedata_signal
			rmm_deb_fee_hk_rd_address_o            => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,             --                                             .rd_address_signal
			rmm_deb_fee_hk_read_o                  => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,                   --                                             .read_signal
			rmm_aeb1_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb1_master_rmap_target.wr_waitrequest_signal
			rmm_aeb1_rmap_target_readdata_i        => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_rmap_target_wr_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb1_rmap_target_write_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb1_rmap_target_writedata_o       => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb1_rmap_target_rd_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb1_rmap_target_read_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb1_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb1_master_fee_hk.wr_waitrequest_signal
			rmm_aeb1_fee_hk_readdata_i             => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_fee_hk_wr_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb1_fee_hk_write_o                => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb1_fee_hk_writedata_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb1_fee_hk_rd_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb1_fee_hk_read_o                 => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb2_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb2_master_rmap_target.wr_waitrequest_signal
			rmm_aeb2_rmap_target_readdata_i        => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_rmap_target_wr_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb2_rmap_target_write_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb2_rmap_target_writedata_o       => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb2_rmap_target_rd_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb2_rmap_target_read_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb2_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb2_master_fee_hk.wr_waitrequest_signal
			rmm_aeb2_fee_hk_readdata_i             => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_fee_hk_wr_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb2_fee_hk_write_o                => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb2_fee_hk_writedata_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb2_fee_hk_rd_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb2_fee_hk_read_o                 => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb3_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb3_master_rmap_target.wr_waitrequest_signal
			rmm_aeb3_rmap_target_readdata_i        => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_rmap_target_wr_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb3_rmap_target_write_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb3_rmap_target_writedata_o       => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb3_rmap_target_rd_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb3_rmap_target_read_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb3_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb3_master_fee_hk.wr_waitrequest_signal
			rmm_aeb3_fee_hk_readdata_i             => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_fee_hk_wr_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb3_fee_hk_write_o                => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb3_fee_hk_writedata_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb3_fee_hk_rd_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb3_fee_hk_read_o                 => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb4_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb4_master_rmap_target.wr_waitrequest_signal
			rmm_aeb4_rmap_target_readdata_i        => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_rmap_target_wr_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb4_rmap_target_write_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb4_rmap_target_writedata_o       => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb4_rmap_target_rd_address_o      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb4_rmap_target_read_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb4_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb4_master_fee_hk.wr_waitrequest_signal
			rmm_aeb4_fee_hk_readdata_i             => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_fee_hk_wr_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb4_fee_hk_write_o                => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb4_fee_hk_writedata_o            => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb4_fee_hk_rd_address_o           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb4_fee_hk_read_o                 => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,                  --                                             .read_signal
			channel_hk_rmap_target_status_o        => communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_status_signal,                 --                   conduit_end_channel_hk_out.rmap_target_status_signal
			channel_hk_rmap_target_indicate_o      => communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_indicate_signal,               --                                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_escape_err_signal,                --                                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_credit_err_signal,                --                                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_parity_err_signal,                --                                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_disconnect_signal,                --                                             .spw_link_disconnect_signal
			channel_hk_spw_link_started_o          => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_started_signal,                   --                                             .spw_link_started_signal
			channel_hk_spw_link_connecting_o       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_connecting_signal,                --                                             .spw_link_connecting_signal
			channel_hk_spw_link_running_o          => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_running_signal,                   --                                             .spw_link_running_signal
			channel_hk_frame_counter_o             => communication_module_v2_ch2_conduit_end_channel_hk_out_frame_counter_signal,                      --                                             .frame_counter_signal
			channel_hk_left_buffer_ccd_number_o    => communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,             --                                             .left_buffer_ccd_number_signal
			channel_hk_right_buffer_ccd_number_o   => communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,            --                                             .right_buffer_ccd_number_signal
			channel_hk_left_buffer_ccd_side_o      => communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,               --                                             .left_buffer_ccd_side_signal
			channel_hk_right_buffer_ccd_side_o     => communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,              --                                             .right_buffer_ccd_side_signal
			channel_hk_err_left_buffer_overflow_o  => communication_module_v2_ch2_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,           --                                             .err_left_buffer_overflow_signal
			channel_hk_err_right_buffer_overflow_o => communication_module_v2_ch2_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,          --                                             .err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_o          => communication_module_v2_ch2_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal,          --             conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
			comm_data_control_data_hold_i          => comm_2_data_control_data_hold_signal,                                                             --                            comm_data_control.data_hold_signal
			comm_measurements_o                    => comm_2_measurements_measurements_signal                                                           --                conduit_end_comm_measurements.measurements_signal
		);

	communication_module_v2_ch3 : component comm_v2_top
		port map (
			reset_sink_reset_i                     => rst_controller_002_reset_out_reset,                                                               --                                   reset_sink.reset
			clock_sink_clk_i                       => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                                   clock_sink.clk
			channel_sync_i                         => comm_3_sync_sync_signal,                                                                          --                     conduit_end_channel_sync.sync_signal
			avs_config_address_i                   => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_address,                     --                       avalon_mm_config_slave.address
			avs_config_write_i                     => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_write,                       --                                             .write
			avs_config_writedata_i                 => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_writedata,                   --                                             .writedata
			avs_config_read_i                      => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_read,                        --                                             .read
			avs_config_readdata_o                  => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_readdata,                    --                                             .readdata
			avs_config_waitrequest_o               => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_waitrequest,                 --                                             .waitrequest
			avm_left_buffer_readdata_i             => communication_module_v2_ch3_avalon_mm_left_buffer_master_readdata,                                --                 avalon_mm_left_buffer_master.readdata
			avm_left_buffer_waitrequest_i          => communication_module_v2_ch3_avalon_mm_left_buffer_master_waitrequest,                             --                                             .waitrequest
			avm_left_buffer_address_o              => communication_module_v2_ch3_avalon_mm_left_buffer_master_address,                                 --                                             .address
			avm_left_buffer_read_o                 => communication_module_v2_ch3_avalon_mm_left_buffer_master_read,                                    --                                             .read
			avm_right_buffer_readdata_i            => communication_module_v2_ch3_avalon_mm_right_buffer_master_readdata,                               --                avalon_mm_right_buffer_master.readdata
			avm_right_buffer_waitrequest_i         => communication_module_v2_ch3_avalon_mm_right_buffer_master_waitrequest,                            --                                             .waitrequest
			avm_right_buffer_address_o             => communication_module_v2_ch3_avalon_mm_right_buffer_master_address,                                --                                             .address
			avm_right_buffer_read_o                => communication_module_v2_ch3_avalon_mm_right_buffer_master_read,                                   --                                             .read
			feeb_interrupt_sender_irq_o            => irq_mapper_receiver3_irq,                                                                         --                        feeb_interrupt_sender.irq
			rmap_interrupt_sender_irq_o            => irq_mapper_receiver12_irq,                                                                        --                        rmap_interrupt_sender.irq
			spw_link_status_started_i              => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --             conduit_end_spacewire_controller.spw_link_status_started_signal
			spw_link_status_connecting_i           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                             .spw_link_status_connecting_signal
			spw_link_status_running_i              => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                             .spw_link_status_running_signal
			spw_link_error_errdisc_i               => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                             .spw_link_error_errdisc_signal
			spw_link_error_errpar_i                => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                             .spw_link_error_errpar_signal
			spw_link_error_erresc_i                => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                             .spw_link_error_erresc_signal
			spw_link_error_errcred_i               => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                             .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_i             => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                             .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_i             => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                             .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_i             => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                             .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_i           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                             .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_i           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                             .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_i            => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                             .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_i            => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                             .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_i             => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                             .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_i           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                             .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_i          => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                             .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_i         => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                             .spw_errinj_ctrl_errinj_ready_signal
			spw_link_command_enable_o              => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --                                             .spw_link_command_enable_signal
			spw_link_command_autostart_o           => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                             .spw_link_command_autostart_signal
			spw_link_command_linkstart_o           => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                             .spw_link_command_linkstart_signal
			spw_link_command_linkdis_o             => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                             .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_o            => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                             .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_o              => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                             .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_o              => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                             .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_o              => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                             .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_o           => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                             .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_o          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                             .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_o           => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                             .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_o           => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                             .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_o         => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                             .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_o         => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                             .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_o          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                             .spw_errinj_ctrl_errinj_code_signal
			rmap_echo_echo_en_o                    => communication_module_v2_ch3_conduit_end_rmap_echo_out_echo_en_signal,                             --                    conduit_end_rmap_echo_out.echo_en_signal
			rmap_echo_echo_id_en_o                 => communication_module_v2_ch3_conduit_end_rmap_echo_out_echo_id_en_signal,                          --                                             .echo_id_en_signal
			rmap_echo_in_fifo_wrflag_o             => communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                      --                                             .in_fifo_wrflag_signal
			rmap_echo_in_fifo_wrdata_o             => communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                      --                                             .in_fifo_wrdata_signal
			rmap_echo_in_fifo_wrreq_o              => communication_module_v2_ch3_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                       --                                             .in_fifo_wrreq_signal
			rmap_echo_out_fifo_wrflag_o            => communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                     --                                             .out_fifo_wrflag_signal
			rmap_echo_out_fifo_wrdata_o            => communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                     --                                             .out_fifo_wrdata_signal
			rmap_echo_out_fifo_wrreq_o             => communication_module_v2_ch3_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                      --                                             .out_fifo_wrreq_signal
			rmm_deb_rmap_target_wr_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                        --  conduit_end_rmap_mem_deb_master_rmap_target.wr_waitrequest_signal
			rmm_deb_rmap_target_readdata_i         => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_rmap_target_rd_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_rmap_target_wr_address_o       => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal,        --                                             .wr_address_signal
			rmm_deb_rmap_target_write_o            => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,             --                                             .write_signal
			rmm_deb_rmap_target_writedata_o        => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,         --                                             .writedata_signal
			rmm_deb_rmap_target_rd_address_o       => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal,        --                                             .rd_address_signal
			rmm_deb_rmap_target_read_o             => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,              --                                             .read_signal
			rmm_deb_fee_hk_wr_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                        --       conduit_end_rmap_mem_deb_master_fee_hk.wr_waitrequest_signal
			rmm_deb_fee_hk_readdata_i              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_fee_hk_rd_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_fee_hk_wr_address_o            => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,             --                                             .wr_address_signal
			rmm_deb_fee_hk_write_o                 => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,                  --                                             .write_signal
			rmm_deb_fee_hk_writedata_o             => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,              --                                             .writedata_signal
			rmm_deb_fee_hk_rd_address_o            => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,             --                                             .rd_address_signal
			rmm_deb_fee_hk_read_o                  => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,                   --                                             .read_signal
			rmm_aeb1_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb1_master_rmap_target.wr_waitrequest_signal
			rmm_aeb1_rmap_target_readdata_i        => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_rmap_target_wr_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb1_rmap_target_write_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb1_rmap_target_writedata_o       => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb1_rmap_target_rd_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb1_rmap_target_read_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb1_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb1_master_fee_hk.wr_waitrequest_signal
			rmm_aeb1_fee_hk_readdata_i             => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_fee_hk_wr_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb1_fee_hk_write_o                => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb1_fee_hk_writedata_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb1_fee_hk_rd_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb1_fee_hk_read_o                 => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb2_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb2_master_rmap_target.wr_waitrequest_signal
			rmm_aeb2_rmap_target_readdata_i        => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_rmap_target_wr_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb2_rmap_target_write_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb2_rmap_target_writedata_o       => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb2_rmap_target_rd_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb2_rmap_target_read_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb2_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb2_master_fee_hk.wr_waitrequest_signal
			rmm_aeb2_fee_hk_readdata_i             => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_fee_hk_wr_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb2_fee_hk_write_o                => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb2_fee_hk_writedata_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb2_fee_hk_rd_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb2_fee_hk_read_o                 => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb3_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb3_master_rmap_target.wr_waitrequest_signal
			rmm_aeb3_rmap_target_readdata_i        => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_rmap_target_wr_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb3_rmap_target_write_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb3_rmap_target_writedata_o       => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb3_rmap_target_rd_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb3_rmap_target_read_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb3_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb3_master_fee_hk.wr_waitrequest_signal
			rmm_aeb3_fee_hk_readdata_i             => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_fee_hk_wr_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb3_fee_hk_write_o                => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb3_fee_hk_writedata_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb3_fee_hk_rd_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb3_fee_hk_read_o                 => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb4_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb4_master_rmap_target.wr_waitrequest_signal
			rmm_aeb4_rmap_target_readdata_i        => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_rmap_target_wr_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb4_rmap_target_write_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb4_rmap_target_writedata_o       => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb4_rmap_target_rd_address_o      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb4_rmap_target_read_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb4_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb4_master_fee_hk.wr_waitrequest_signal
			rmm_aeb4_fee_hk_readdata_i             => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_fee_hk_wr_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb4_fee_hk_write_o                => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb4_fee_hk_writedata_o            => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb4_fee_hk_rd_address_o           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb4_fee_hk_read_o                 => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,                  --                                             .read_signal
			channel_hk_rmap_target_status_o        => communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_status_signal,                 --                   conduit_end_channel_hk_out.rmap_target_status_signal
			channel_hk_rmap_target_indicate_o      => communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_indicate_signal,               --                                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_escape_err_signal,                --                                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_credit_err_signal,                --                                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_parity_err_signal,                --                                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_disconnect_signal,                --                                             .spw_link_disconnect_signal
			channel_hk_spw_link_started_o          => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_started_signal,                   --                                             .spw_link_started_signal
			channel_hk_spw_link_connecting_o       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_connecting_signal,                --                                             .spw_link_connecting_signal
			channel_hk_spw_link_running_o          => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_running_signal,                   --                                             .spw_link_running_signal
			channel_hk_frame_counter_o             => communication_module_v2_ch3_conduit_end_channel_hk_out_frame_counter_signal,                      --                                             .frame_counter_signal
			channel_hk_left_buffer_ccd_number_o    => communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,             --                                             .left_buffer_ccd_number_signal
			channel_hk_right_buffer_ccd_number_o   => communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,            --                                             .right_buffer_ccd_number_signal
			channel_hk_left_buffer_ccd_side_o      => communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,               --                                             .left_buffer_ccd_side_signal
			channel_hk_right_buffer_ccd_side_o     => communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,              --                                             .right_buffer_ccd_side_signal
			channel_hk_err_left_buffer_overflow_o  => communication_module_v2_ch3_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,           --                                             .err_left_buffer_overflow_signal
			channel_hk_err_right_buffer_overflow_o => communication_module_v2_ch3_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,          --                                             .err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_o          => communication_module_v2_ch3_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal,          --             conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
			comm_data_control_data_hold_i          => comm_3_data_control_data_hold_signal,                                                             --                            comm_data_control.data_hold_signal
			comm_measurements_o                    => comm_3_measurements_measurements_signal                                                           --                conduit_end_comm_measurements.measurements_signal
		);

	communication_module_v2_ch4 : component comm_v2_top
		port map (
			reset_sink_reset_i                     => rst_controller_002_reset_out_reset,                                                               --                                   reset_sink.reset
			clock_sink_clk_i                       => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                                   clock_sink.clk
			channel_sync_i                         => comm_4_sync_sync_signal,                                                                          --                     conduit_end_channel_sync.sync_signal
			avs_config_address_i                   => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_address,                     --                       avalon_mm_config_slave.address
			avs_config_write_i                     => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_write,                       --                                             .write
			avs_config_writedata_i                 => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_writedata,                   --                                             .writedata
			avs_config_read_i                      => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_read,                        --                                             .read
			avs_config_readdata_o                  => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_readdata,                    --                                             .readdata
			avs_config_waitrequest_o               => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_waitrequest,                 --                                             .waitrequest
			avm_left_buffer_readdata_i             => communication_module_v2_ch4_avalon_mm_left_buffer_master_readdata,                                --                 avalon_mm_left_buffer_master.readdata
			avm_left_buffer_waitrequest_i          => communication_module_v2_ch4_avalon_mm_left_buffer_master_waitrequest,                             --                                             .waitrequest
			avm_left_buffer_address_o              => communication_module_v2_ch4_avalon_mm_left_buffer_master_address,                                 --                                             .address
			avm_left_buffer_read_o                 => communication_module_v2_ch4_avalon_mm_left_buffer_master_read,                                    --                                             .read
			avm_right_buffer_readdata_i            => communication_module_v2_ch4_avalon_mm_right_buffer_master_readdata,                               --                avalon_mm_right_buffer_master.readdata
			avm_right_buffer_waitrequest_i         => communication_module_v2_ch4_avalon_mm_right_buffer_master_waitrequest,                            --                                             .waitrequest
			avm_right_buffer_address_o             => communication_module_v2_ch4_avalon_mm_right_buffer_master_address,                                --                                             .address
			avm_right_buffer_read_o                => communication_module_v2_ch4_avalon_mm_right_buffer_master_read,                                   --                                             .read
			feeb_interrupt_sender_irq_o            => irq_mapper_receiver2_irq,                                                                         --                        feeb_interrupt_sender.irq
			rmap_interrupt_sender_irq_o            => irq_mapper_receiver11_irq,                                                                        --                        rmap_interrupt_sender.irq
			spw_link_status_started_i              => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --             conduit_end_spacewire_controller.spw_link_status_started_signal
			spw_link_status_connecting_i           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                             .spw_link_status_connecting_signal
			spw_link_status_running_i              => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                             .spw_link_status_running_signal
			spw_link_error_errdisc_i               => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                             .spw_link_error_errdisc_signal
			spw_link_error_errpar_i                => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                             .spw_link_error_errpar_signal
			spw_link_error_erresc_i                => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                             .spw_link_error_erresc_signal
			spw_link_error_errcred_i               => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                             .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_i             => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                             .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_i             => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                             .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_i             => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                             .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_i           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                             .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_i           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                             .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_i            => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                             .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_i            => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                             .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_i             => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                             .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_i           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                             .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_i          => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                             .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_i         => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                             .spw_errinj_ctrl_errinj_ready_signal
			spw_link_command_enable_o              => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --                                             .spw_link_command_enable_signal
			spw_link_command_autostart_o           => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                             .spw_link_command_autostart_signal
			spw_link_command_linkstart_o           => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                             .spw_link_command_linkstart_signal
			spw_link_command_linkdis_o             => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                             .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_o            => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                             .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_o              => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                             .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_o              => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                             .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_o              => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                             .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_o           => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                             .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_o          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                             .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_o           => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                             .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_o           => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                             .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_o         => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                             .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_o         => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                             .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_o          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                             .spw_errinj_ctrl_errinj_code_signal
			rmap_echo_echo_en_o                    => communication_module_v2_ch4_conduit_end_rmap_echo_out_echo_en_signal,                             --                    conduit_end_rmap_echo_out.echo_en_signal
			rmap_echo_echo_id_en_o                 => communication_module_v2_ch4_conduit_end_rmap_echo_out_echo_id_en_signal,                          --                                             .echo_id_en_signal
			rmap_echo_in_fifo_wrflag_o             => communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrflag_signal,                      --                                             .in_fifo_wrflag_signal
			rmap_echo_in_fifo_wrdata_o             => communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrdata_signal,                      --                                             .in_fifo_wrdata_signal
			rmap_echo_in_fifo_wrreq_o              => communication_module_v2_ch4_conduit_end_rmap_echo_out_in_fifo_wrreq_signal,                       --                                             .in_fifo_wrreq_signal
			rmap_echo_out_fifo_wrflag_o            => communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrflag_signal,                     --                                             .out_fifo_wrflag_signal
			rmap_echo_out_fifo_wrdata_o            => communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrdata_signal,                     --                                             .out_fifo_wrdata_signal
			rmap_echo_out_fifo_wrreq_o             => communication_module_v2_ch4_conduit_end_rmap_echo_out_out_fifo_wrreq_signal,                      --                                             .out_fifo_wrreq_signal
			rmm_deb_rmap_target_wr_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                        --  conduit_end_rmap_mem_deb_master_rmap_target.wr_waitrequest_signal
			rmm_deb_rmap_target_readdata_i         => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_rmap_target_rd_waitrequest_i   => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_rmap_target_wr_address_o       => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal,        --                                             .wr_address_signal
			rmm_deb_rmap_target_write_o            => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,             --                                             .write_signal
			rmm_deb_rmap_target_writedata_o        => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,         --                                             .writedata_signal
			rmm_deb_rmap_target_rd_address_o       => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal,        --                                             .rd_address_signal
			rmm_deb_rmap_target_read_o             => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,              --                                             .read_signal
			rmm_deb_fee_hk_wr_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                        --       conduit_end_rmap_mem_deb_master_fee_hk.wr_waitrequest_signal
			rmm_deb_fee_hk_readdata_i              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_readdata_signal,                              --                                             .readdata_signal
			rmm_deb_fee_hk_rd_waitrequest_i        => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                        --                                             .rd_waitrequest_signal
			rmm_deb_fee_hk_wr_address_o            => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,             --                                             .wr_address_signal
			rmm_deb_fee_hk_write_o                 => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,                  --                                             .write_signal
			rmm_deb_fee_hk_writedata_o             => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,              --                                             .writedata_signal
			rmm_deb_fee_hk_rd_address_o            => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,             --                                             .rd_address_signal
			rmm_deb_fee_hk_read_o                  => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,                   --                                             .read_signal
			rmm_aeb1_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb1_master_rmap_target.wr_waitrequest_signal
			rmm_aeb1_rmap_target_readdata_i        => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_rmap_target_wr_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb1_rmap_target_write_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb1_rmap_target_writedata_o       => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb1_rmap_target_rd_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb1_rmap_target_read_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb1_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb1_master_fee_hk.wr_waitrequest_signal
			rmm_aeb1_fee_hk_readdata_i             => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb1_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb1_fee_hk_wr_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb1_fee_hk_write_o                => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb1_fee_hk_writedata_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb1_fee_hk_rd_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb1_fee_hk_read_o                 => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb2_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb2_master_rmap_target.wr_waitrequest_signal
			rmm_aeb2_rmap_target_readdata_i        => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_rmap_target_wr_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb2_rmap_target_write_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb2_rmap_target_writedata_o       => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb2_rmap_target_rd_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb2_rmap_target_read_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb2_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb2_master_fee_hk.wr_waitrequest_signal
			rmm_aeb2_fee_hk_readdata_i             => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb2_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb2_fee_hk_wr_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb2_fee_hk_write_o                => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb2_fee_hk_writedata_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb2_fee_hk_rd_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb2_fee_hk_read_o                 => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb3_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb3_master_rmap_target.wr_waitrequest_signal
			rmm_aeb3_rmap_target_readdata_i        => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_rmap_target_wr_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb3_rmap_target_write_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb3_rmap_target_writedata_o       => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb3_rmap_target_rd_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb3_rmap_target_read_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb3_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb3_master_fee_hk.wr_waitrequest_signal
			rmm_aeb3_fee_hk_readdata_i             => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb3_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb3_fee_hk_wr_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb3_fee_hk_write_o                => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb3_fee_hk_writedata_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb3_fee_hk_rd_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb3_fee_hk_read_o                 => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,                  --                                             .read_signal
			rmm_aeb4_rmap_target_wr_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                      -- conduit_end_rmap_mem_aeb4_master_rmap_target.wr_waitrequest_signal
			rmm_aeb4_rmap_target_readdata_i        => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_rmap_target_rd_waitrequest_i  => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_rmap_target_wr_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal,       --                                             .wr_address_signal
			rmm_aeb4_rmap_target_write_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,            --                                             .write_signal
			rmm_aeb4_rmap_target_writedata_o       => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,        --                                             .writedata_signal
			rmm_aeb4_rmap_target_rd_address_o      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal,       --                                             .rd_address_signal
			rmm_aeb4_rmap_target_read_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,             --                                             .read_signal
			rmm_aeb4_fee_hk_wr_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                      --      conduit_end_rmap_mem_aeb4_master_fee_hk.wr_waitrequest_signal
			rmm_aeb4_fee_hk_readdata_i             => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_readdata_signal,                            --                                             .readdata_signal
			rmm_aeb4_fee_hk_rd_waitrequest_i       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                      --                                             .rd_waitrequest_signal
			rmm_aeb4_fee_hk_wr_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,            --                                             .wr_address_signal
			rmm_aeb4_fee_hk_write_o                => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,                 --                                             .write_signal
			rmm_aeb4_fee_hk_writedata_o            => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,             --                                             .writedata_signal
			rmm_aeb4_fee_hk_rd_address_o           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,            --                                             .rd_address_signal
			rmm_aeb4_fee_hk_read_o                 => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,                  --                                             .read_signal
			channel_hk_rmap_target_status_o        => communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_status_signal,                 --                   conduit_end_channel_hk_out.rmap_target_status_signal
			channel_hk_rmap_target_indicate_o      => communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_indicate_signal,               --                                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_escape_err_signal,                --                                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_credit_err_signal,                --                                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_parity_err_signal,                --                                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_disconnect_signal,                --                                             .spw_link_disconnect_signal
			channel_hk_spw_link_started_o          => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_started_signal,                   --                                             .spw_link_started_signal
			channel_hk_spw_link_connecting_o       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_connecting_signal,                --                                             .spw_link_connecting_signal
			channel_hk_spw_link_running_o          => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_running_signal,                   --                                             .spw_link_running_signal
			channel_hk_frame_counter_o             => communication_module_v2_ch4_conduit_end_channel_hk_out_frame_counter_signal,                      --                                             .frame_counter_signal
			channel_hk_left_buffer_ccd_number_o    => communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,             --                                             .left_buffer_ccd_number_signal
			channel_hk_right_buffer_ccd_number_o   => communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,            --                                             .right_buffer_ccd_number_signal
			channel_hk_left_buffer_ccd_side_o      => communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,               --                                             .left_buffer_ccd_side_signal
			channel_hk_right_buffer_ccd_side_o     => communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,              --                                             .right_buffer_ccd_side_signal
			channel_hk_err_left_buffer_overflow_o  => communication_module_v2_ch4_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,           --                                             .err_left_buffer_overflow_signal
			channel_hk_err_right_buffer_overflow_o => communication_module_v2_ch4_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,          --                                             .err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_o          => communication_module_v2_ch4_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal,          --             conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
			comm_data_control_data_hold_i          => comm_4_data_control_data_hold_signal,                                                             --                            comm_data_control.data_hold_signal
			comm_measurements_o                    => comm_4_measurements_measurements_signal                                                           --                conduit_end_comm_measurements.measurements_signal
		);

	ftdi_umft601a_module : component ftdi_usb3_top
		port map (
			clock_sink_clk_i                      => m2_ddr2_memory_afi_half_clk_clk,                                        --              clock_sink.clk
			reset_sink_reset_i                    => rst_controller_002_reset_out_reset,                                     --              reset_sink.reset
			umft601a_clock_sink_clk_i             => ftdi_clk_clk,                                                           --     umft601a_clock_sink.clk
			umft601a_clock_pin_i                  => umft601a_pins_umft_clock_signal,                                        --   conduit_umft601a_pins.umft_clock_signal
			umft601a_txe_n_pin_i                  => umft601a_pins_umft_txe_n_signal,                                        --                        .umft_txe_n_signal
			umft601a_rxf_n_pin_i                  => umft601a_pins_umft_rxf_n_signal,                                        --                        .umft_rxf_n_signal
			umft601a_data_bus_io                  => umft601a_pins_umft_data_signal,                                         --                        .umft_data_signal
			umft601a_be_bus_io                    => umft601a_pins_umft_be_signal,                                           --                        .umft_be_signal
			umft601a_wakeup_n_pin_io              => umft601a_pins_umft_wakeup_n_signal,                                     --                        .umft_wakeup_n_signal
			umft601a_gpio_bus_io                  => umft601a_pins_umft_gpio_bus_signal,                                     --                        .umft_gpio_bus_signal
			umft601a_reset_n_pin_o                => umft601a_pins_umft_reset_n_signal,                                      --                        .umft_reset_n_signal
			umft601a_wr_n_pin_o                   => umft601a_pins_umft_wr_n_signal,                                         --                        .umft_wr_n_signal
			umft601a_rd_n_pin_o                   => umft601a_pins_umft_rd_n_signal,                                         --                        .umft_rd_n_signal
			umft601a_oe_n_pin_o                   => umft601a_pins_umft_oe_n_signal,                                         --                        .umft_oe_n_signal
			umft601a_siwu_n_pin_o                 => umft601a_pins_umft_siwu_n_signal,                                       --                        .umft_siwu_n_signal
			avalon_slave_config_address_i         => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_address,     --     avalon_slave_config.address
			avalon_slave_config_write_i           => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_write,       --                        .write
			avalon_slave_config_writedata_i       => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_writedata,   --                        .writedata
			avalon_slave_config_read_i            => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_read,        --                        .read
			avalon_slave_config_readdata_o        => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_readdata,    --                        .readdata
			avalon_slave_config_waitrequest_o     => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_waitrequest, --                        .waitrequest
			avalon_master_data_readdata_i         => ftdi_umft601a_module_avalon_master_data_readdata,                       --      avalon_master_data.readdata
			avalon_master_data_waitrequest_i      => ftdi_umft601a_module_avalon_master_data_waitrequest,                    --                        .waitrequest
			avalon_master_data_address_o          => ftdi_umft601a_module_avalon_master_data_address,                        --                        .address
			avalon_master_data_read_o             => ftdi_umft601a_module_avalon_master_data_read,                           --                        .read
			avalon_master_data_write_o            => ftdi_umft601a_module_avalon_master_data_write,                          --                        .write
			avalon_master_data_writedata_o        => ftdi_umft601a_module_avalon_master_data_writedata,                      --                        .writedata
			avalon_imgt_master_data_waitrequest_i => ftdi_umft601a_module_avalon_imgt_master_data_waitrequest,               -- avalon_imgt_master_data.waitrequest
			avalon_imgt_master_data_address_o     => ftdi_umft601a_module_avalon_imgt_master_data_address,                   --                        .address
			avalon_imgt_master_data_write_o       => ftdi_umft601a_module_avalon_imgt_master_data_write,                     --                        .write
			avalon_imgt_master_data_writedata_o   => ftdi_umft601a_module_avalon_imgt_master_data_writedata,                 --                        .writedata
			rx_interrupt_sender_irq_o             => irq_mapper_receiver13_irq,                                              --     rx_interrupt_sender.irq
			tx_interrupt_sender_irq_o             => irq_mapper_receiver15_irq,                                              --     tx_interrupt_sender.irq
			ftdi_data_control_sync_pulse_i        => ftdi_data_control_sync_pulse_signal,                                    --       ftdi_data_control.sync_pulse_signal
			ftdi_data_control_data_hold_o         => ftdi_data_control_data_hold_signal                                      --                        .data_hold_signal
		);

	memory_filler : component mfil_memory_filler_top
		port map (
			clock_sink_clk_i                  => m2_ddr2_memory_afi_half_clk_clk,                                 --          clock_sink.clk
			reset_sink_reset_i                => rst_controller_002_reset_out_reset,                              --          reset_sink.reset
			avalon_slave_config_address_i     => mm_interconnect_1_memory_filler_avalon_slave_config_address,     -- avalon_slave_config.address
			avalon_slave_config_byteenable_i  => mm_interconnect_1_memory_filler_avalon_slave_config_byteenable,  --                    .byteenable
			avalon_slave_config_write_i       => mm_interconnect_1_memory_filler_avalon_slave_config_write,       --                    .write
			avalon_slave_config_writedata_i   => mm_interconnect_1_memory_filler_avalon_slave_config_writedata,   --                    .writedata
			avalon_slave_config_read_i        => mm_interconnect_1_memory_filler_avalon_slave_config_read,        --                    .read
			avalon_slave_config_readdata_o    => mm_interconnect_1_memory_filler_avalon_slave_config_readdata,    --                    .readdata
			avalon_slave_config_waitrequest_o => mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest, --                    .waitrequest
			avalon_master_data_waitrequest_i  => memory_filler_avalon_master_data_waitrequest,                    --  avalon_master_data.waitrequest
			avalon_master_data_address_o      => memory_filler_avalon_master_data_address,                        --                    .address
			avalon_master_data_write_o        => memory_filler_avalon_master_data_write,                          --                    .write
			avalon_master_data_writedata_o    => memory_filler_avalon_master_data_writedata                       --                    .writedata
		);

	spacewire_channel_a : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_a_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_a_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_a_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_a_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_a_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_a_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_a_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_a_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_a_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_a_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_a_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_a_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_b : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_b_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_b_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_b_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_b_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_b_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_b_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_b_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_b_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_b_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_b_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_b_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_b_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_c : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_c_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_c_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_c_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_c_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_c_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_c_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_c_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_c_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_c_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_c_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_c_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_c_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_d : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_d_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_d_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_d_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_d_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_d_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_d_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_d_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_d_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_d_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_d_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_d_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_d_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_e : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_e_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_e_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_e_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_e_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_e_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_e_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_e_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_e_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_e_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_e_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_e_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_e_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_f : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_f_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_f_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_f_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_f_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_f_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_f_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_f_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_f_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_f_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_f_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_f_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_f_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_g : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_g_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_g_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_g_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_g_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_g_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_g_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_g_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_g_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_g_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_g_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_g_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_g_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_channel_h : component spwc_spacewire_channel_top
		port map (
			reset_i                        => rst_controller_003_reset_out_reset,                                                         --                    reset_sink.reset
			clk_100_i                      => m2_ddr2_memory_afi_half_clk_clk,                                                            --             clock_sink_100mhz.clk
			clk_200_i                      => m2_ddr2_memory_afi_clk_clk,                                                                 --             clock_sink_200mhz.clk
			spw_lvds_p_data_in_i           => spwc_h_lvds_spw_lvds_p_data_in_signal,                                                      --    conduit_end_spacewire_lvds.spw_lvds_p_data_in_signal
			spw_lvds_n_data_in_i           => spwc_h_lvds_spw_lvds_n_data_in_signal,                                                      --                              .spw_lvds_n_data_in_signal
			spw_lvds_p_data_out_o          => spwc_h_lvds_spw_lvds_p_data_out_signal,                                                     --                              .spw_lvds_p_data_out_signal
			spw_lvds_n_data_out_o          => spwc_h_lvds_spw_lvds_n_data_out_signal,                                                     --                              .spw_lvds_n_data_out_signal
			spw_lvds_p_strobe_out_o        => spwc_h_lvds_spw_lvds_p_strobe_out_signal,                                                   --                              .spw_lvds_p_strobe_out_signal
			spw_lvds_n_strobe_out_o        => spwc_h_lvds_spw_lvds_n_strobe_out_signal,                                                   --                              .spw_lvds_n_strobe_out_signal
			spw_lvds_p_strobe_in_i         => spwc_h_lvds_spw_lvds_p_strobe_in_signal,                                                    --                              .spw_lvds_p_strobe_in_signal
			spw_lvds_n_strobe_in_i         => spwc_h_lvds_spw_lvds_n_strobe_in_signal,                                                    --                              .spw_lvds_n_strobe_in_signal
			spw_rx_enable_i                => spwc_h_enable_spw_rx_enable_signal,                                                         --  conduit_end_spacewire_enable.spw_rx_enable_signal
			spw_tx_enable_i                => spwc_h_enable_spw_tx_enable_signal,                                                         --                              .spw_tx_enable_signal
			spw_red_status_led_o           => spwc_h_leds_spw_red_status_led_signal,                                                      --    conduit_end_spacewire_leds.spw_red_status_led_signal
			spw_green_status_led_o         => spwc_h_leds_spw_green_status_led_signal,                                                    --                              .spw_green_status_led_signal
			spw_link_command_enable_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,      -- conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,   --                              .spw_link_command_autostart_signal
			spw_link_command_linkstart_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,   --                              .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i     => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,     --                              .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i    => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,    --                              .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,      --                              .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,      --                              .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,      --                              .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,   --                              .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i  => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,  --                              .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,   --                              .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,   --                              .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal, --                              .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal, --                              .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i  => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal,  --                              .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o      => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal,           --                              .spw_link_status_started_signal
			spw_link_status_connecting_o   => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal,        --                              .spw_link_status_connecting_signal
			spw_link_status_running_o      => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal,           --                              .spw_link_status_running_signal
			spw_link_error_errdisc_o       => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,            --                              .spw_link_error_errdisc_signal
			spw_link_error_errpar_o        => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal,             --                              .spw_link_error_errpar_signal
			spw_link_error_erresc_o        => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal,             --                              .spw_link_error_erresc_signal
			spw_link_error_errcred_o       => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal,            --                              .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,          --                              .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,          --                              .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,          --                              .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,        --                              .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,        --                              .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o    => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,         --                              .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o    => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,         --                              .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o     => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,          --                              .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,        --                              .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o  => spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,       --                              .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o => spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal       --                              .spw_errinj_ctrl_errinj_ready_signal
		);

	spacewire_demux_ch1 : component spwd_spacewire_demux_top
		port map (
			reset_i                            => rst_controller_002_reset_out_reset,                                                               --                         reset_sink.reset
			clock_i                            => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                         clock_sink.clk
			demux_select_i                     => spwd_ch1_select_demux_select_signal,                                                              --           conduit_end_demux_select.demux_select_signal
			spw_link_command_enable_i          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --      conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i       => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                   .spw_link_command_autostart_signal
			spw_link_command_linkstart_i       => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                   .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i         => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                   .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i        => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                   .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                   .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                   .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i          => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                   .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i       => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                   .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i      => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                   .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i       => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                   .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i       => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                   .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i     => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i     => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i      => communication_module_v2_ch1_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o          => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --                                   .spw_link_status_started_signal
			spw_link_status_connecting_o       => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_link_status_running_o          => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_link_error_errdisc_o           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_link_error_errpar_o            => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_link_error_erresc_o            => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_link_error_errcred_o           => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o         => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o         => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o         => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o       => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o       => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o        => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o        => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o         => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o       => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o      => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o     => spacewire_demux_ch1_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_status_started_i      => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_0.spw_link_status_started_signal
			spw_ct0_link_status_connecting_i   => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct0_link_status_running_i      => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct0_link_error_errdisc_i       => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct0_link_error_errpar_i        => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct0_link_error_erresc_i        => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct0_link_error_errcred_i       => spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct0_timecode_rx_tick_out_i     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct0_timecode_rx_ctrl_out_i     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct0_timecode_rx_time_out_i     => spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct0_data_rx_status_rxvalid_i   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct0_data_rx_status_rxhalff_i   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct0_data_rx_status_rxflag_i    => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct0_data_rx_status_rxdata_i    => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct0_data_tx_status_txrdy_i     => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct0_data_tx_status_txhalff_i   => spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct0_errinj_ctrl_errinj_busy_i  => spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct0_errinj_ctrl_errinj_ready_i => spacewire_channel_a_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_command_enable_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct0_link_command_autostart_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct0_link_command_linkstart_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct0_link_command_linkdis_o     => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct0_link_command_txdivcnt_o    => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct0_timecode_tx_tick_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct0_timecode_tx_ctrl_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct0_timecode_tx_time_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct0_data_rx_command_rxread_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct0_data_tx_command_txwrite_o  => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct0_data_tx_command_txflag_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct0_data_tx_command_txdata_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct0_errinj_ctrl_start_errinj_o => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct0_errinj_ctrl_reset_errinj_o => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct0_errinj_ctrl_errinj_code_o  => spacewire_demux_ch1_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,        --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_ct1_link_status_started_i      => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_1.spw_link_status_started_signal
			spw_ct1_link_status_connecting_i   => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct1_link_status_running_i      => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct1_link_error_errdisc_i       => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct1_link_error_errpar_i        => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct1_link_error_erresc_i        => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct1_link_error_errcred_i       => spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct1_timecode_rx_tick_out_i     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct1_timecode_rx_ctrl_out_i     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct1_timecode_rx_time_out_i     => spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct1_data_rx_status_rxvalid_i   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct1_data_rx_status_rxhalff_i   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct1_data_rx_status_rxflag_i    => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct1_data_rx_status_rxdata_i    => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct1_data_tx_status_txrdy_i     => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct1_data_tx_status_txhalff_i   => spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct1_errinj_ctrl_errinj_busy_i  => spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct1_errinj_ctrl_errinj_ready_i => spacewire_channel_e_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct1_link_command_enable_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct1_link_command_autostart_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct1_link_command_linkstart_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct1_link_command_linkdis_o     => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct1_link_command_txdivcnt_o    => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct1_timecode_tx_tick_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct1_timecode_tx_ctrl_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct1_timecode_tx_time_in_o      => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct1_data_rx_command_rxread_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct1_data_tx_command_txwrite_o  => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct1_data_tx_command_txflag_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct1_data_tx_command_txdata_o   => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct1_errinj_ctrl_start_errinj_o => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct1_errinj_ctrl_reset_errinj_o => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct1_errinj_ctrl_errinj_code_o  => spacewire_demux_ch1_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal         --                                   .spw_errinj_ctrl_errinj_code_signal
		);

	spacewire_demux_ch2 : component spwd_spacewire_demux_top
		port map (
			reset_i                            => rst_controller_002_reset_out_reset,                                                               --                         reset_sink.reset
			clock_i                            => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                         clock_sink.clk
			demux_select_i                     => spwd_ch2_select_demux_select_signal,                                                              --           conduit_end_demux_select.demux_select_signal
			spw_link_command_enable_i          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --      conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i       => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                   .spw_link_command_autostart_signal
			spw_link_command_linkstart_i       => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                   .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i         => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                   .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i        => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                   .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                   .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                   .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i          => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                   .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i       => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                   .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i      => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                   .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i       => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                   .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i       => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                   .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i     => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i     => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i      => communication_module_v2_ch2_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o          => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --                                   .spw_link_status_started_signal
			spw_link_status_connecting_o       => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_link_status_running_o          => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_link_error_errdisc_o           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_link_error_errpar_o            => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_link_error_erresc_o            => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_link_error_errcred_o           => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o         => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o         => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o         => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o       => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o       => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o        => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o        => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o         => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o       => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o      => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o     => spacewire_demux_ch2_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_status_started_i      => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_0.spw_link_status_started_signal
			spw_ct0_link_status_connecting_i   => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct0_link_status_running_i      => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct0_link_error_errdisc_i       => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct0_link_error_errpar_i        => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct0_link_error_erresc_i        => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct0_link_error_errcred_i       => spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct0_timecode_rx_tick_out_i     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct0_timecode_rx_ctrl_out_i     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct0_timecode_rx_time_out_i     => spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct0_data_rx_status_rxvalid_i   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct0_data_rx_status_rxhalff_i   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct0_data_rx_status_rxflag_i    => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct0_data_rx_status_rxdata_i    => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct0_data_tx_status_txrdy_i     => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct0_data_tx_status_txhalff_i   => spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct0_errinj_ctrl_errinj_busy_i  => spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct0_errinj_ctrl_errinj_ready_i => spacewire_channel_b_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_command_enable_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct0_link_command_autostart_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct0_link_command_linkstart_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct0_link_command_linkdis_o     => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct0_link_command_txdivcnt_o    => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct0_timecode_tx_tick_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct0_timecode_tx_ctrl_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct0_timecode_tx_time_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct0_data_rx_command_rxread_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct0_data_tx_command_txwrite_o  => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct0_data_tx_command_txflag_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct0_data_tx_command_txdata_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct0_errinj_ctrl_start_errinj_o => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct0_errinj_ctrl_reset_errinj_o => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct0_errinj_ctrl_errinj_code_o  => spacewire_demux_ch2_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,        --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_ct1_link_status_started_i      => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_1.spw_link_status_started_signal
			spw_ct1_link_status_connecting_i   => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct1_link_status_running_i      => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct1_link_error_errdisc_i       => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct1_link_error_errpar_i        => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct1_link_error_erresc_i        => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct1_link_error_errcred_i       => spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct1_timecode_rx_tick_out_i     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct1_timecode_rx_ctrl_out_i     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct1_timecode_rx_time_out_i     => spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct1_data_rx_status_rxvalid_i   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct1_data_rx_status_rxhalff_i   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct1_data_rx_status_rxflag_i    => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct1_data_rx_status_rxdata_i    => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct1_data_tx_status_txrdy_i     => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct1_data_tx_status_txhalff_i   => spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct1_errinj_ctrl_errinj_busy_i  => spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct1_errinj_ctrl_errinj_ready_i => spacewire_channel_f_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct1_link_command_enable_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct1_link_command_autostart_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct1_link_command_linkstart_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct1_link_command_linkdis_o     => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct1_link_command_txdivcnt_o    => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct1_timecode_tx_tick_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct1_timecode_tx_ctrl_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct1_timecode_tx_time_in_o      => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct1_data_rx_command_rxread_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct1_data_tx_command_txwrite_o  => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct1_data_tx_command_txflag_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct1_data_tx_command_txdata_o   => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct1_errinj_ctrl_start_errinj_o => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct1_errinj_ctrl_reset_errinj_o => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct1_errinj_ctrl_errinj_code_o  => spacewire_demux_ch2_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal         --                                   .spw_errinj_ctrl_errinj_code_signal
		);

	spacewire_demux_ch3 : component spwd_spacewire_demux_top
		port map (
			reset_i                            => rst_controller_002_reset_out_reset,                                                               --                         reset_sink.reset
			clock_i                            => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                         clock_sink.clk
			demux_select_i                     => spwd_ch3_select_demux_select_signal,                                                              --           conduit_end_demux_select.demux_select_signal
			spw_link_command_enable_i          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --      conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i       => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                   .spw_link_command_autostart_signal
			spw_link_command_linkstart_i       => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                   .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i         => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                   .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i        => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                   .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                   .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                   .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i          => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                   .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i       => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                   .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i      => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                   .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i       => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                   .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i       => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                   .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i     => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i     => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i      => communication_module_v2_ch3_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o          => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --                                   .spw_link_status_started_signal
			spw_link_status_connecting_o       => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_link_status_running_o          => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_link_error_errdisc_o           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_link_error_errpar_o            => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_link_error_erresc_o            => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_link_error_errcred_o           => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o         => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o         => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o         => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o       => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o       => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o        => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o        => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o         => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o       => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o      => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o     => spacewire_demux_ch3_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_status_started_i      => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_0.spw_link_status_started_signal
			spw_ct0_link_status_connecting_i   => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct0_link_status_running_i      => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct0_link_error_errdisc_i       => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct0_link_error_errpar_i        => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct0_link_error_erresc_i        => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct0_link_error_errcred_i       => spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct0_timecode_rx_tick_out_i     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct0_timecode_rx_ctrl_out_i     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct0_timecode_rx_time_out_i     => spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct0_data_rx_status_rxvalid_i   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct0_data_rx_status_rxhalff_i   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct0_data_rx_status_rxflag_i    => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct0_data_rx_status_rxdata_i    => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct0_data_tx_status_txrdy_i     => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct0_data_tx_status_txhalff_i   => spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct0_errinj_ctrl_errinj_busy_i  => spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct0_errinj_ctrl_errinj_ready_i => spacewire_channel_c_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_command_enable_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct0_link_command_autostart_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct0_link_command_linkstart_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct0_link_command_linkdis_o     => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct0_link_command_txdivcnt_o    => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct0_timecode_tx_tick_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct0_timecode_tx_ctrl_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct0_timecode_tx_time_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct0_data_rx_command_rxread_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct0_data_tx_command_txwrite_o  => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct0_data_tx_command_txflag_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct0_data_tx_command_txdata_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct0_errinj_ctrl_start_errinj_o => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct0_errinj_ctrl_reset_errinj_o => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct0_errinj_ctrl_errinj_code_o  => spacewire_demux_ch3_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,        --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_ct1_link_status_started_i      => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_1.spw_link_status_started_signal
			spw_ct1_link_status_connecting_i   => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct1_link_status_running_i      => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct1_link_error_errdisc_i       => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct1_link_error_errpar_i        => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct1_link_error_erresc_i        => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct1_link_error_errcred_i       => spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct1_timecode_rx_tick_out_i     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct1_timecode_rx_ctrl_out_i     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct1_timecode_rx_time_out_i     => spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct1_data_rx_status_rxvalid_i   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct1_data_rx_status_rxhalff_i   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct1_data_rx_status_rxflag_i    => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct1_data_rx_status_rxdata_i    => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct1_data_tx_status_txrdy_i     => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct1_data_tx_status_txhalff_i   => spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct1_errinj_ctrl_errinj_busy_i  => spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct1_errinj_ctrl_errinj_ready_i => spacewire_channel_g_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct1_link_command_enable_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct1_link_command_autostart_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct1_link_command_linkstart_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct1_link_command_linkdis_o     => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct1_link_command_txdivcnt_o    => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct1_timecode_tx_tick_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct1_timecode_tx_ctrl_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct1_timecode_tx_time_in_o      => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct1_data_rx_command_rxread_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct1_data_tx_command_txwrite_o  => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct1_data_tx_command_txflag_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct1_data_tx_command_txdata_o   => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct1_errinj_ctrl_start_errinj_o => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct1_errinj_ctrl_reset_errinj_o => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct1_errinj_ctrl_errinj_code_o  => spacewire_demux_ch3_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal         --                                   .spw_errinj_ctrl_errinj_code_signal
		);

	spacewire_demux_ch4 : component spwd_spacewire_demux_top
		port map (
			reset_i                            => rst_controller_002_reset_out_reset,                                                               --                         reset_sink.reset
			clock_i                            => m2_ddr2_memory_afi_half_clk_clk,                                                                  --                         clock_sink.clk
			demux_select_i                     => spwd_ch4_select_demux_select_signal,                                                              --           conduit_end_demux_select.demux_select_signal
			spw_link_command_enable_i          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_enable_signal,      --      conduit_end_spacewire_channel.spw_link_command_enable_signal
			spw_link_command_autostart_i       => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_autostart_signal,   --                                   .spw_link_command_autostart_signal
			spw_link_command_linkstart_i       => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal,   --                                   .spw_link_command_linkstart_signal
			spw_link_command_linkdis_i         => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal,     --                                   .spw_link_command_linkdis_signal
			spw_link_command_txdivcnt_i        => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal,    --                                   .spw_link_command_txdivcnt_signal
			spw_timecode_tx_tick_in_i          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal,      --                                   .spw_timecode_tx_tick_in_signal
			spw_timecode_tx_ctrl_in_i          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal,      --                                   .spw_timecode_tx_ctrl_in_signal
			spw_timecode_tx_time_in_i          => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal,      --                                   .spw_timecode_tx_time_in_signal
			spw_data_rx_command_rxread_i       => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal,   --                                   .spw_data_rx_command_rxread_signal
			spw_data_tx_command_txwrite_i      => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal,  --                                   .spw_data_tx_command_txwrite_signal
			spw_data_tx_command_txflag_i       => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal,   --                                   .spw_data_tx_command_txflag_signal
			spw_data_tx_command_txdata_i       => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal,   --                                   .spw_data_tx_command_txdata_signal
			spw_errinj_ctrl_start_errinj_i     => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_start_errinj_signal, --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_errinj_ctrl_reset_errinj_i     => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_reset_errinj_signal, --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_errinj_ctrl_errinj_code_i      => communication_module_v2_ch4_conduit_end_spacewire_controller_spw_errinj_ctrl_errinj_code_signal,  --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_link_status_started_o          => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_started_signal,                 --                                   .spw_link_status_started_signal
			spw_link_status_connecting_o       => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_link_status_running_o          => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_link_error_errdisc_o           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_link_error_errpar_o            => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_link_error_erresc_o            => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_link_error_errcred_o           => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_timecode_rx_tick_out_o         => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_timecode_rx_ctrl_out_o         => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_timecode_rx_time_out_o         => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_data_rx_status_rxvalid_o       => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_data_rx_status_rxhalff_o       => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_data_rx_status_rxflag_o        => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_data_rx_status_rxdata_o        => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_data_tx_status_txrdy_o         => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_data_tx_status_txhalff_o       => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_errinj_ctrl_errinj_busy_o      => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_errinj_ctrl_errinj_ready_o     => spacewire_demux_ch4_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_status_started_i      => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_0.spw_link_status_started_signal
			spw_ct0_link_status_connecting_i   => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct0_link_status_running_i      => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct0_link_error_errdisc_i       => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct0_link_error_errpar_i        => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct0_link_error_erresc_i        => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct0_link_error_errcred_i       => spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct0_timecode_rx_tick_out_i     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct0_timecode_rx_ctrl_out_i     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct0_timecode_rx_time_out_i     => spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct0_data_rx_status_rxvalid_i   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct0_data_rx_status_rxhalff_i   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct0_data_rx_status_rxflag_i    => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct0_data_rx_status_rxdata_i    => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct0_data_tx_status_txrdy_i     => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct0_data_tx_status_txhalff_i   => spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct0_errinj_ctrl_errinj_busy_i  => spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct0_errinj_ctrl_errinj_ready_i => spacewire_channel_d_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct0_link_command_enable_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct0_link_command_autostart_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct0_link_command_linkstart_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct0_link_command_linkdis_o     => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct0_link_command_txdivcnt_o    => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct0_timecode_tx_tick_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct0_timecode_tx_ctrl_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct0_timecode_tx_time_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct0_data_rx_command_rxread_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct0_data_tx_command_txwrite_o  => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct0_data_tx_command_txflag_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct0_data_tx_command_txdata_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct0_errinj_ctrl_start_errinj_o => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct0_errinj_ctrl_reset_errinj_o => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct0_errinj_ctrl_errinj_code_o  => spacewire_demux_ch4_conduit_end_spacewire_controller_0_spw_errinj_ctrl_errinj_code_signal,        --                                   .spw_errinj_ctrl_errinj_code_signal
			spw_ct1_link_status_started_i      => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal,                 -- conduit_end_spacewire_controller_1.spw_link_status_started_signal
			spw_ct1_link_status_connecting_i   => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal,              --                                   .spw_link_status_connecting_signal
			spw_ct1_link_status_running_i      => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal,                 --                                   .spw_link_status_running_signal
			spw_ct1_link_error_errdisc_i       => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal,                  --                                   .spw_link_error_errdisc_signal
			spw_ct1_link_error_errpar_i        => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal,                   --                                   .spw_link_error_errpar_signal
			spw_ct1_link_error_erresc_i        => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal,                   --                                   .spw_link_error_erresc_signal
			spw_ct1_link_error_errcred_i       => spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal,                  --                                   .spw_link_error_errcred_signal
			spw_ct1_timecode_rx_tick_out_i     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal,                --                                   .spw_timecode_rx_tick_out_signal
			spw_ct1_timecode_rx_ctrl_out_i     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal,                --                                   .spw_timecode_rx_ctrl_out_signal
			spw_ct1_timecode_rx_time_out_i     => spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal,                --                                   .spw_timecode_rx_time_out_signal
			spw_ct1_data_rx_status_rxvalid_i   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal,              --                                   .spw_data_rx_status_rxvalid_signal
			spw_ct1_data_rx_status_rxhalff_i   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal,              --                                   .spw_data_rx_status_rxhalff_signal
			spw_ct1_data_rx_status_rxflag_i    => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal,               --                                   .spw_data_rx_status_rxflag_signal
			spw_ct1_data_rx_status_rxdata_i    => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal,               --                                   .spw_data_rx_status_rxdata_signal
			spw_ct1_data_tx_status_txrdy_i     => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal,                --                                   .spw_data_tx_status_txrdy_signal
			spw_ct1_data_tx_status_txhalff_i   => spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal,              --                                   .spw_data_tx_status_txhalff_signal
			spw_ct1_errinj_ctrl_errinj_busy_i  => spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_busy_signal,             --                                   .spw_errinj_ctrl_errinj_busy_signal
			spw_ct1_errinj_ctrl_errinj_ready_i => spacewire_channel_h_conduit_end_spacewire_channel_spw_errinj_ctrl_errinj_ready_signal,            --                                   .spw_errinj_ctrl_errinj_ready_signal
			spw_ct1_link_command_enable_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_enable_signal,            --                                   .spw_link_command_enable_signal
			spw_ct1_link_command_autostart_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_autostart_signal,         --                                   .spw_link_command_autostart_signal
			spw_ct1_link_command_linkstart_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkstart_signal,         --                                   .spw_link_command_linkstart_signal
			spw_ct1_link_command_linkdis_o     => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_linkdis_signal,           --                                   .spw_link_command_linkdis_signal
			spw_ct1_link_command_txdivcnt_o    => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_link_command_txdivcnt_signal,          --                                   .spw_link_command_txdivcnt_signal
			spw_ct1_timecode_tx_tick_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_tick_in_signal,            --                                   .spw_timecode_tx_tick_in_signal
			spw_ct1_timecode_tx_ctrl_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_ctrl_in_signal,            --                                   .spw_timecode_tx_ctrl_in_signal
			spw_ct1_timecode_tx_time_in_o      => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_timecode_tx_time_in_signal,            --                                   .spw_timecode_tx_time_in_signal
			spw_ct1_data_rx_command_rxread_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_rx_command_rxread_signal,         --                                   .spw_data_rx_command_rxread_signal
			spw_ct1_data_tx_command_txwrite_o  => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txwrite_signal,        --                                   .spw_data_tx_command_txwrite_signal
			spw_ct1_data_tx_command_txflag_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txflag_signal,         --                                   .spw_data_tx_command_txflag_signal
			spw_ct1_data_tx_command_txdata_o   => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_data_tx_command_txdata_signal,         --                                   .spw_data_tx_command_txdata_signal
			spw_ct1_errinj_ctrl_start_errinj_o => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_start_errinj_signal,       --                                   .spw_errinj_ctrl_start_errinj_signal
			spw_ct1_errinj_ctrl_reset_errinj_o => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_reset_errinj_signal,       --                                   .spw_errinj_ctrl_reset_errinj_signal
			spw_ct1_errinj_ctrl_errinj_code_o  => spacewire_demux_ch4_conduit_end_spacewire_controller_1_spw_errinj_ctrl_errinj_code_signal         --                                   .spw_errinj_ctrl_errinj_code_signal
		);

	clock_bridge_afi_50 : component mebx_qsys_project_clock_bridge_afi_50
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk50_clk,                                              --   m0_clk.clk
			m0_reset         => rst_controller_001_reset_out_reset,                     -- m0_reset.reset
			s0_clk           => m2_ddr2_memory_afi_half_clk_clk,                        --   s0_clk.clk
			s0_reset         => rst_controller_002_reset_out_reset,                     -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_1_clock_bridge_afi_50_s0_address,       --         .address
			s0_write         => mm_interconnect_1_clock_bridge_afi_50_s0_write,         --         .write
			s0_read          => mm_interconnect_1_clock_bridge_afi_50_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => clock_bridge_afi_50_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => clock_bridge_afi_50_m0_readdata,                        --         .readdata
			m0_readdatavalid => clock_bridge_afi_50_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => clock_bridge_afi_50_m0_burstcount,                      --         .burstcount
			m0_writedata     => clock_bridge_afi_50_m0_writedata,                       --         .writedata
			m0_address       => clock_bridge_afi_50_m0_address,                         --         .address
			m0_write         => clock_bridge_afi_50_m0_write,                           --         .write
			m0_read          => clock_bridge_afi_50_m0_read,                            --         .read
			m0_byteenable    => clock_bridge_afi_50_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => clock_bridge_afi_50_m0_debugaccess                      --         .debugaccess
		);

	csense_adc_fo : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                          --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_2_csense_adc_fo_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_adc_fo_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_adc_fo_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_adc_fo_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_adc_fo_s1_readdata,        --                    .readdata
			out_port   => csense_adc_fo_export                                -- external_connection.export
		);

	csense_cs_n : component MebX_Qsys_Project_csense_cs_n
		port map (
			clk        => clk50_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_2_csense_cs_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_cs_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_cs_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_cs_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_cs_n_s1_readdata,        --                    .readdata
			out_port   => csense_cs_n_export                                -- external_connection.export
		);

	csense_sck : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sck_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sck_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sck_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sck_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sck_s1_readdata,        --                    .readdata
			out_port   => csense_sck_export                                -- external_connection.export
		);

	csense_sdi : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sdi_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sdi_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sdi_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sdi_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sdi_s1_readdata,        --                    .readdata
			out_port   => csense_sdi_export                                -- external_connection.export
		);

	csense_sdo : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_csense_sdo_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_csense_sdo_s1_readdata,     --                    .readdata
			in_port  => csense_sdo_export                             -- external_connection.export
		);

	ddr2_address_span_extender : component altera_address_span_extender
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 29,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 8,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			clk                  => m2_ddr2_memory_afi_half_clk_clk,                                           --           clock.clk
			reset                => rst_controller_002_reset_out_reset,                                        --           reset.reset
			avs_s0_address       => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => ddr2_address_span_extender_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => ddr2_address_span_extender_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => ddr2_address_span_extender_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => ddr2_address_span_extender_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => ddr2_address_span_extender_expanded_master_write,                          --                .write
			avm_m0_writedata     => ddr2_address_span_extender_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => ddr2_address_span_extender_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => ddr2_address_span_extender_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => ddr2_address_span_extender_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_read        => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                    --            cntl.read
			avs_cntl_readdata    => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                --                .readdata
			avs_cntl_write       => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                   --                .write
			avs_cntl_writedata   => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,               --                .writedata
			avs_cntl_byteenable  => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,              --                .byteenable
			avs_cntl_address     => "0"                                                                        --     (terminated)
		);

	ext_flash : component MebX_Qsys_Project_ext_flash
		generic map (
			TCM_ADDRESS_W                  => 26,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 100,
			TCM_WRITE_WAIT                 => 100,
			TCM_SETUP_WAIT                 => 25,
			TCM_DATA_HOLD                  => 20,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => m2_ddr2_memory_afi_half_clk_clk,               --   clk.clk
			reset_reset          => rst_controller_004_reset_out_reset,            -- reset.reset
			uas_address          => mm_interconnect_1_ext_flash_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_1_ext_flash_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_1_ext_flash_uas_read,          --      .read
			uas_write            => mm_interconnect_1_ext_flash_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_1_ext_flash_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_1_ext_flash_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_1_ext_flash_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_1_ext_flash_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_1_ext_flash_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_1_ext_flash_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_1_ext_flash_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ext_flash_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_n_out       => ext_flash_tcm_read_n_out,                      --      .read_n_out
			tcm_chipselect_n_out => ext_flash_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ext_flash_tcm_request,                         --      .request
			tcm_grant            => ext_flash_tcm_grant,                           --      .grant
			tcm_address_out      => ext_flash_tcm_address_out,                     --      .address_out
			tcm_data_out         => ext_flash_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ext_flash_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ext_flash_tcm_data_in                          --      .data_in
		);

	jtag_uart_0 : component MebX_Qsys_Project_jtag_uart_0
		port map (
			clk            => m2_ddr2_memory_afi_half_clk_clk,                                 --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver4_irq                                         --               irq.irq
		);

	m1_clock_bridge : component mebx_qsys_project_m1_clock_bridge
		generic map (
			DATA_WIDTH          => 256,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 31,
			BURSTCOUNT_WIDTH    => 3,
			COMMAND_FIFO_DEPTH  => 8,
			RESPONSE_FIFO_DEPTH => 8,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => m1_ddr2_memory_afi_half_clk_clk,                    --   m0_clk.clk
			m0_reset         => rst_controller_005_reset_out_reset,                 -- m0_reset.reset
			s0_clk           => m2_ddr2_memory_afi_half_clk_clk,                    --   s0_clk.clk
			s0_reset         => rst_controller_002_reset_out_reset,                 -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_m1_clock_bridge_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_m1_clock_bridge_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_m1_clock_bridge_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_m1_clock_bridge_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_m1_clock_bridge_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_m1_clock_bridge_s0_address,       --         .address
			s0_write         => mm_interconnect_0_m1_clock_bridge_s0_write,         --         .write
			s0_read          => mm_interconnect_0_m1_clock_bridge_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_m1_clock_bridge_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_m1_clock_bridge_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => m1_clock_bridge_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => m1_clock_bridge_m0_readdata,                        --         .readdata
			m0_readdatavalid => m1_clock_bridge_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => m1_clock_bridge_m0_burstcount,                      --         .burstcount
			m0_writedata     => m1_clock_bridge_m0_writedata,                       --         .writedata
			m0_address       => m1_clock_bridge_m0_address,                         --         .address
			m0_write         => m1_clock_bridge_m0_write,                           --         .write
			m0_read          => m1_clock_bridge_m0_read,                            --         .read
			m0_byteenable    => m1_clock_bridge_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => m1_clock_bridge_m0_debugaccess                      --         .debugaccess
		);

	m1_ddr2_i2c_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m1_ddr2_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => m1_ddr2_i2c_scl_export                                -- external_connection.export
		);

	m1_ddr2_i2c_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m1_ddr2_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => m1_ddr2_i2c_sda_export                                -- external_connection.export
		);

	m1_ddr2_memory : component MebX_Qsys_Project_m1_ddr2_memory
		port map (
			pll_ref_clk        => m1_ddr2_memory_pll_ref_clk_clk,                          --      pll_ref_clk.clk
			global_reset_n     => rst_reset_n,                                             --     global_reset.reset_n
			soft_reset_n       => rst_reset_n,                                             --       soft_reset.reset_n
			afi_clk            => m1_ddr2_memory_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk       => m1_ddr2_memory_afi_half_clk_clk,                         --     afi_half_clk.clk
			afi_reset_n        => open,                                                    --        afi_reset.reset_n
			afi_reset_export_n => open,                                                    -- afi_reset_export.reset_n
			mem_a              => m1_ddr2_memory_mem_a,                                    --           memory.mem_a
			mem_ba             => m1_ddr2_memory_mem_ba,                                   --                 .mem_ba
			mem_ck             => m1_ddr2_memory_mem_ck,                                   --                 .mem_ck
			mem_ck_n           => m1_ddr2_memory_mem_ck_n,                                 --                 .mem_ck_n
			mem_cke            => m1_ddr2_memory_mem_cke,                                  --                 .mem_cke
			mem_cs_n           => m1_ddr2_memory_mem_cs_n,                                 --                 .mem_cs_n
			mem_dm             => m1_ddr2_memory_mem_dm,                                   --                 .mem_dm
			mem_ras_n          => m1_ddr2_memory_mem_ras_n,                                --                 .mem_ras_n
			mem_cas_n          => m1_ddr2_memory_mem_cas_n,                                --                 .mem_cas_n
			mem_we_n           => m1_ddr2_memory_mem_we_n,                                 --                 .mem_we_n
			mem_dq             => m1_ddr2_memory_mem_dq,                                   --                 .mem_dq
			mem_dqs            => m1_ddr2_memory_mem_dqs,                                  --                 .mem_dqs
			mem_dqs_n          => m1_ddr2_memory_mem_dqs_n,                                --                 .mem_dqs_n
			mem_odt            => m1_ddr2_memory_mem_odt,                                  --                 .mem_odt
			avl_ready          => m1_ddr2_memory_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin     => mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr           => mm_interconnect_3_m1_ddr2_memory_avl_address,            --                 .address
			avl_rdata_valid    => mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata          => mm_interconnect_3_m1_ddr2_memory_avl_readdata,           --                 .readdata
			avl_wdata          => mm_interconnect_3_m1_ddr2_memory_avl_writedata,          --                 .writedata
			avl_be             => mm_interconnect_3_m1_ddr2_memory_avl_byteenable,         --                 .byteenable
			avl_read_req       => mm_interconnect_3_m1_ddr2_memory_avl_read,               --                 .read
			avl_write_req      => mm_interconnect_3_m1_ddr2_memory_avl_write,              --                 .write
			avl_size           => mm_interconnect_3_m1_ddr2_memory_avl_burstcount,         --                 .burstcount
			local_init_done    => m1_ddr2_memory_status_local_init_done,                   --           status.local_init_done
			local_cal_success  => m1_ddr2_memory_status_local_cal_success,                 --                 .local_cal_success
			local_cal_fail     => m1_ddr2_memory_status_local_cal_fail,                    --                 .local_cal_fail
			oct_rdn            => m1_ddr2_oct_rdn,                                         --              oct.rdn
			oct_rup            => m1_ddr2_oct_rup                                          --                 .rup
		);

	m2_ddr2_i2c_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m2_ddr2_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => m2_ddr2_i2c_scl_export                                -- external_connection.export
		);

	m2_ddr2_i2c_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m2_ddr2_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => m2_ddr2_i2c_sda_export                                -- external_connection.export
		);

	m2_ddr2_memory : component MebX_Qsys_Project_m2_ddr2_memory
		port map (
			pll_ref_clk               => clk50_clk,                                               --      pll_ref_clk.clk
			global_reset_n            => rst_reset_n,                                             --     global_reset.reset_n
			soft_reset_n              => rst_reset_n,                                             --       soft_reset.reset_n
			afi_clk                   => m2_ddr2_memory_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk              => m2_ddr2_memory_afi_half_clk_clk,                         --     afi_half_clk.clk
			afi_reset_n               => open,                                                    --        afi_reset.reset_n
			afi_reset_export_n        => open,                                                    -- afi_reset_export.reset_n
			mem_a                     => m2_ddr2_memory_mem_a,                                    --           memory.mem_a
			mem_ba                    => m2_ddr2_memory_mem_ba,                                   --                 .mem_ba
			mem_ck                    => m2_ddr2_memory_mem_ck,                                   --                 .mem_ck
			mem_ck_n                  => m2_ddr2_memory_mem_ck_n,                                 --                 .mem_ck_n
			mem_cke                   => m2_ddr2_memory_mem_cke,                                  --                 .mem_cke
			mem_cs_n                  => m2_ddr2_memory_mem_cs_n,                                 --                 .mem_cs_n
			mem_dm                    => m2_ddr2_memory_mem_dm,                                   --                 .mem_dm
			mem_ras_n                 => m2_ddr2_memory_mem_ras_n,                                --                 .mem_ras_n
			mem_cas_n                 => m2_ddr2_memory_mem_cas_n,                                --                 .mem_cas_n
			mem_we_n                  => m2_ddr2_memory_mem_we_n,                                 --                 .mem_we_n
			mem_dq                    => m2_ddr2_memory_mem_dq,                                   --                 .mem_dq
			mem_dqs                   => m2_ddr2_memory_mem_dqs,                                  --                 .mem_dqs
			mem_dqs_n                 => m2_ddr2_memory_mem_dqs_n,                                --                 .mem_dqs_n
			mem_odt                   => m2_ddr2_memory_mem_odt,                                  --                 .mem_odt
			avl_ready                 => m2_ddr2_memory_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin            => mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr                  => mm_interconnect_0_m2_ddr2_memory_avl_address,            --                 .address
			avl_rdata_valid           => mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata                 => mm_interconnect_0_m2_ddr2_memory_avl_readdata,           --                 .readdata
			avl_wdata                 => mm_interconnect_0_m2_ddr2_memory_avl_writedata,          --                 .writedata
			avl_be                    => mm_interconnect_0_m2_ddr2_memory_avl_byteenable,         --                 .byteenable
			avl_read_req              => mm_interconnect_0_m2_ddr2_memory_avl_read,               --                 .read
			avl_write_req             => mm_interconnect_0_m2_ddr2_memory_avl_write,              --                 .write
			avl_size                  => mm_interconnect_0_m2_ddr2_memory_avl_burstcount,         --                 .burstcount
			local_init_done           => m2_ddr2_memory_status_local_init_done,                   --           status.local_init_done
			local_cal_success         => m2_ddr2_memory_status_local_cal_success,                 --                 .local_cal_success
			local_cal_fail            => m2_ddr2_memory_status_local_cal_fail,                    --                 .local_cal_fail
			oct_rdn                   => m2_ddr2_oct_rdn,                                         --              oct.rdn
			oct_rup                   => m2_ddr2_oct_rup,                                         --                 .rup
			pll_mem_clk               => m2_ddr2_memory_pll_sharing_pll_mem_clk,                  --      pll_sharing.pll_mem_clk
			pll_write_clk             => m2_ddr2_memory_pll_sharing_pll_write_clk,                --                 .pll_write_clk
			pll_locked                => m2_ddr2_memory_pll_sharing_pll_locked,                   --                 .pll_locked
			pll_write_clk_pre_phy_clk => m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk,    --                 .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          => m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,             --                 .pll_addr_cmd_clk
			pll_avl_clk               => m2_ddr2_memory_pll_sharing_pll_avl_clk,                  --                 .pll_avl_clk
			pll_config_clk            => m2_ddr2_memory_pll_sharing_pll_config_clk,               --                 .pll_config_clk
			dll_pll_locked            => m2_ddr2_memory_dll_sharing_dll_pll_locked,               --      dll_sharing.dll_pll_locked
			dll_delayctrl             => m2_ddr2_memory_dll_sharing_dll_delayctrl                 --                 .dll_delayctrl
		);

	nios2_gen2_0 : component MebX_Qsys_Project_nios2_gen2_0
		port map (
			clk                                 => m2_ddr2_memory_afi_half_clk_clk,                            --                       clk.clk
			reset_n                             => rst_controller_006_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_006_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_burstcount                        => nios2_gen2_0_instruction_master_burstcount,                 --                          .burstcount
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory : component MebX_Qsys_Project_onchip_memory
		port map (
			clk        => m2_ddr2_memory_afi_half_clk_clk,               --   clk1.clk
			address    => mm_interconnect_1_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_1_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_1_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_002_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_002_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	pio_button : component MebX_Qsys_Project_pio_BUTTON
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_button_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_pio_button_s1_readdata,     --                    .readdata
			in_port  => button_export                                 -- external_connection.export
		);

	pio_dip : component MebX_Qsys_Project_pio_DIP
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_dip_s1_address,         --                  s1.address
			readdata => mm_interconnect_2_pio_dip_s1_readdata,        --                    .readdata
			in_port  => dip_export                                    -- external_connection.export
		);

	pio_ext : component MebX_Qsys_Project_pio_EXT
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_ext_s1_address,         --                  s1.address
			readdata => mm_interconnect_2_pio_ext_s1_readdata,        --                    .readdata
			in_port  => ext_export                                    -- external_connection.export
		);

	pio_led : component MebX_Qsys_Project_pio_LED
		port map (
			clk        => clk50_clk,                                    --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_led_s1_readdata,        --                    .readdata
			out_port   => led_de4_export                                -- external_connection.export
		);

	pio_led_painel : component MebX_Qsys_Project_pio_LED_painel
		port map (
			clk        => clk50_clk,                                           --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_2_pio_led_painel_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_led_painel_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_led_painel_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_led_painel_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_led_painel_s1_readdata,        --                    .readdata
			out_port   => led_painel_export                                    -- external_connection.export
		);

	pio_ctrl_io_lvds : component MebX_Qsys_Project_pio_ctrl_io_lvds
		port map (
			clk        => clk50_clk,                                             --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_2_pio_ctrl_io_lvds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata,        --                    .readdata
			out_port   => ctrl_io_lvds_export                                    -- external_connection.export
		);

	pio_ftdi_umft601a_module_reset : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                                           --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_readdata,        --                    .readdata
			out_port   => pio_ftdi_umft601a_module_reset_export                                -- external_connection.export
		);

	pio_iso_logic_signal_enable : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => mm_interconnect_2_pio_iso_logic_signal_enable_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_iso_logic_signal_enable_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_iso_logic_signal_enable_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_iso_logic_signal_enable_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_iso_logic_signal_enable_s1_readdata,        --                    .readdata
			out_port   => pio_iso_logic_signal_enable_export                                -- external_connection.export
		);

	pio_spw_demux_ch_1_select : component MebX_Qsys_Project_pio_spw_demux_ch_1_select
		port map (
			clk        => clk50_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_readdata,        --                    .readdata
			out_port   => pio_spw_demux_ch_1_select_export                                -- external_connection.export
		);

	pio_spw_demux_ch_2_select : component MebX_Qsys_Project_pio_spw_demux_ch_1_select
		port map (
			clk        => clk50_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_readdata,        --                    .readdata
			out_port   => pio_spw_demux_ch_2_select_export                                -- external_connection.export
		);

	pio_spw_demux_ch_3_select : component MebX_Qsys_Project_pio_spw_demux_ch_1_select
		port map (
			clk        => clk50_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_readdata,        --                    .readdata
			out_port   => pio_spw_demux_ch_3_select_export                                -- external_connection.export
		);

	pio_spw_demux_ch_4_select : component MebX_Qsys_Project_pio_spw_demux_ch_1_select
		port map (
			clk        => clk50_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_readdata,        --                    .readdata
			out_port   => pio_spw_demux_ch_4_select_export                                -- external_connection.export
		);

	rmap_mem_ffee_aeb_1_area : component farm_rmap_memory_ffee_aeb_area_top
		port map (
			reset_i                     => rst_controller_002_reset_out_reset,                                                         --                   reset_sink.reset
			clk_100_i                   => m2_ddr2_memory_afi_half_clk_clk,                                                            --            clock_sink_100mhz.clk
			avs_rmap_0_address_i        => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address,                     --          avalon_rmap_slave_0.address
			avs_rmap_0_write_i          => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write,                       --                             .write
			avs_rmap_0_read_i           => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read,                        --                             .read
			avs_rmap_0_readdata_o       => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata,                    --                             .readdata
			avs_rmap_0_writedata_i      => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata,                   --                             .writedata
			avs_rmap_0_waitrequest_o    => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest,                 --                             .waitrequest
			rms_rmap_0_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_0.wr_address_signal
			rms_rmap_0_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_0_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_0_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_0_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_0_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_0_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_readdata_signal,                      --                             .readdata_signal
			rms_rmap_0_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_1_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_1.wr_address_signal
			rms_rmap_1_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_1_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_1_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_1_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_1_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_1_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_readdata_signal,                      --                             .readdata_signal
			rms_rmap_1_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_2_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_2.wr_address_signal
			rms_rmap_2_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_2_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_2_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_2_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_2_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_2_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_readdata_signal,                      --                             .readdata_signal
			rms_rmap_2_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_3_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_3.wr_address_signal
			rms_rmap_3_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_3_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_3_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_3_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_3_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_3_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_readdata_signal,                      --                             .readdata_signal
			rms_rmap_3_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_4_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_4.wr_address_signal
			rms_rmap_4_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_4_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_4_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_4_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_4_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_4_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_readdata_signal,                      --                             .readdata_signal
			rms_rmap_4_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_5_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_5.wr_address_signal
			rms_rmap_5_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_5_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_5_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_5_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_5_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_5_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_readdata_signal,                      --                             .readdata_signal
			rms_rmap_5_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_6_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_6.wr_address_signal
			rms_rmap_6_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_6_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_6_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_6_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_6_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_6_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_readdata_signal,                      --                             .readdata_signal
			rms_rmap_6_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_7_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_7.wr_address_signal
			rms_rmap_7_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_7_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_7_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_7_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb1_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_7_wr_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_7_readdata_o       => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_readdata_signal,                      --                             .readdata_signal
			rms_rmap_7_rd_waitrequest_o => rmap_mem_ffee_aeb_1_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                 --                             .rd_waitrequest_signal
		);

	rmap_mem_ffee_aeb_2_area : component farm_rmap_memory_ffee_aeb_area_top
		port map (
			reset_i                     => rst_controller_002_reset_out_reset,                                                         --                   reset_sink.reset
			clk_100_i                   => m2_ddr2_memory_afi_half_clk_clk,                                                            --            clock_sink_100mhz.clk
			avs_rmap_0_address_i        => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address,                     --          avalon_rmap_slave_0.address
			avs_rmap_0_write_i          => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write,                       --                             .write
			avs_rmap_0_read_i           => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read,                        --                             .read
			avs_rmap_0_readdata_o       => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata,                    --                             .readdata
			avs_rmap_0_writedata_i      => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata,                   --                             .writedata
			avs_rmap_0_waitrequest_o    => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest,                 --                             .waitrequest
			rms_rmap_0_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_0.wr_address_signal
			rms_rmap_0_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_0_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_0_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_0_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_0_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_0_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_readdata_signal,                      --                             .readdata_signal
			rms_rmap_0_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_1_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_1.wr_address_signal
			rms_rmap_1_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_1_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_1_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_1_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_1_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_1_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_readdata_signal,                      --                             .readdata_signal
			rms_rmap_1_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_2_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_2.wr_address_signal
			rms_rmap_2_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_2_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_2_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_2_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_2_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_2_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_readdata_signal,                      --                             .readdata_signal
			rms_rmap_2_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_3_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_3.wr_address_signal
			rms_rmap_3_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_3_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_3_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_3_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_3_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_3_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_readdata_signal,                      --                             .readdata_signal
			rms_rmap_3_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_4_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_4.wr_address_signal
			rms_rmap_4_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_4_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_4_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_4_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_4_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_4_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_readdata_signal,                      --                             .readdata_signal
			rms_rmap_4_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_5_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_5.wr_address_signal
			rms_rmap_5_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_5_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_5_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_5_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_5_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_5_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_readdata_signal,                      --                             .readdata_signal
			rms_rmap_5_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_6_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_6.wr_address_signal
			rms_rmap_6_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_6_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_6_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_6_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_6_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_6_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_readdata_signal,                      --                             .readdata_signal
			rms_rmap_6_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_7_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_7.wr_address_signal
			rms_rmap_7_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_7_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_7_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_7_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb2_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_7_wr_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_7_readdata_o       => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_readdata_signal,                      --                             .readdata_signal
			rms_rmap_7_rd_waitrequest_o => rmap_mem_ffee_aeb_2_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                 --                             .rd_waitrequest_signal
		);

	rmap_mem_ffee_aeb_3_area : component farm_rmap_memory_ffee_aeb_area_top
		port map (
			reset_i                     => rst_controller_002_reset_out_reset,                                                         --                   reset_sink.reset
			clk_100_i                   => m2_ddr2_memory_afi_half_clk_clk,                                                            --            clock_sink_100mhz.clk
			avs_rmap_0_address_i        => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address,                     --          avalon_rmap_slave_0.address
			avs_rmap_0_write_i          => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write,                       --                             .write
			avs_rmap_0_read_i           => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read,                        --                             .read
			avs_rmap_0_readdata_o       => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata,                    --                             .readdata
			avs_rmap_0_writedata_i      => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata,                   --                             .writedata
			avs_rmap_0_waitrequest_o    => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest,                 --                             .waitrequest
			rms_rmap_0_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_0.wr_address_signal
			rms_rmap_0_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_0_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_0_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_0_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_0_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_0_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_readdata_signal,                      --                             .readdata_signal
			rms_rmap_0_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_1_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_1.wr_address_signal
			rms_rmap_1_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_1_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_1_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_1_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_1_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_1_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_readdata_signal,                      --                             .readdata_signal
			rms_rmap_1_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_2_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_2.wr_address_signal
			rms_rmap_2_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_2_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_2_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_2_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_2_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_2_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_readdata_signal,                      --                             .readdata_signal
			rms_rmap_2_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_3_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_3.wr_address_signal
			rms_rmap_3_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_3_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_3_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_3_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_3_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_3_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_readdata_signal,                      --                             .readdata_signal
			rms_rmap_3_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_4_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_4.wr_address_signal
			rms_rmap_4_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_4_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_4_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_4_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_4_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_4_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_readdata_signal,                      --                             .readdata_signal
			rms_rmap_4_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_5_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_5.wr_address_signal
			rms_rmap_5_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_5_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_5_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_5_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_5_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_5_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_readdata_signal,                      --                             .readdata_signal
			rms_rmap_5_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_6_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_6.wr_address_signal
			rms_rmap_6_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_6_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_6_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_6_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_6_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_6_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_readdata_signal,                      --                             .readdata_signal
			rms_rmap_6_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_7_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_7.wr_address_signal
			rms_rmap_7_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_7_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_7_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_7_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb3_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_7_wr_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_7_readdata_o       => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_readdata_signal,                      --                             .readdata_signal
			rms_rmap_7_rd_waitrequest_o => rmap_mem_ffee_aeb_3_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                 --                             .rd_waitrequest_signal
		);

	rmap_mem_ffee_aeb_4_area : component farm_rmap_memory_ffee_aeb_area_top
		port map (
			reset_i                     => rst_controller_002_reset_out_reset,                                                         --                   reset_sink.reset
			clk_100_i                   => m2_ddr2_memory_afi_half_clk_clk,                                                            --            clock_sink_100mhz.clk
			avs_rmap_0_address_i        => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address,                     --          avalon_rmap_slave_0.address
			avs_rmap_0_write_i          => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write,                       --                             .write
			avs_rmap_0_read_i           => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read,                        --                             .read
			avs_rmap_0_readdata_o       => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata,                    --                             .readdata
			avs_rmap_0_writedata_i      => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata,                   --                             .writedata
			avs_rmap_0_waitrequest_o    => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest,                 --                             .waitrequest
			rms_rmap_0_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_0.wr_address_signal
			rms_rmap_0_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_0_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_0_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_0_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_0_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_0_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_readdata_signal,                      --                             .readdata_signal
			rms_rmap_0_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_1_wr_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_1.wr_address_signal
			rms_rmap_1_write_i          => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_1_writedata_i      => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_1_rd_address_i     => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_1_read_i           => communication_module_v2_ch1_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_1_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_1_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_readdata_signal,                      --                             .readdata_signal
			rms_rmap_1_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_2_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_2.wr_address_signal
			rms_rmap_2_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_2_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_2_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_2_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_2_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_2_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_readdata_signal,                      --                             .readdata_signal
			rms_rmap_2_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_3_wr_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_3.wr_address_signal
			rms_rmap_3_write_i          => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_3_writedata_i      => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_3_rd_address_i     => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_3_read_i           => communication_module_v2_ch2_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_3_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_3_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_readdata_signal,                      --                             .readdata_signal
			rms_rmap_3_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_4_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_4.wr_address_signal
			rms_rmap_4_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_4_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_4_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_4_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_4_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_4_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_readdata_signal,                      --                             .readdata_signal
			rms_rmap_4_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_5_wr_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_5.wr_address_signal
			rms_rmap_5_write_i          => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_5_writedata_i      => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_5_rd_address_i     => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_5_read_i           => communication_module_v2_ch3_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_5_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_5_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_readdata_signal,                      --                             .readdata_signal
			rms_rmap_5_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_6_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_wr_address_signal, -- conduit_end_rmap_mem_slave_6.wr_address_signal
			rms_rmap_6_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_write_signal,      --                             .write_signal
			rms_rmap_6_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_writedata_signal,  --                             .writedata_signal
			rms_rmap_6_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_rd_address_signal, --                             .rd_address_signal
			rms_rmap_6_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_rmap_target_read_signal,       --                             .read_signal
			rms_rmap_6_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_6_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_readdata_signal,                      --                             .readdata_signal
			rms_rmap_6_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                --                             .rd_waitrequest_signal
			rms_rmap_7_wr_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_wr_address_signal,      -- conduit_end_rmap_mem_slave_7.wr_address_signal
			rms_rmap_7_write_i          => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_write_signal,           --                             .write_signal
			rms_rmap_7_writedata_i      => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_writedata_signal,       --                             .writedata_signal
			rms_rmap_7_rd_address_i     => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_rd_address_signal,      --                             .rd_address_signal
			rms_rmap_7_read_i           => communication_module_v2_ch4_conduit_end_rmap_mem_aeb4_master_fee_hk_read_signal,            --                             .read_signal
			rms_rmap_7_wr_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                --                             .wr_waitrequest_signal
			rms_rmap_7_readdata_o       => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_readdata_signal,                      --                             .readdata_signal
			rms_rmap_7_rd_waitrequest_o => rmap_mem_ffee_aeb_4_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal                 --                             .rd_waitrequest_signal
		);

	rmap_mem_ffee_deb_area : component fdrm_rmap_memory_ffee_deb_area_top
		port map (
			reset_i                                  => rst_controller_002_reset_out_reset,                                                        --                      reset_sink.reset
			clk_100_i                                => m2_ddr2_memory_afi_half_clk_clk,                                                           --               clock_sink_100mhz.clk
			avs_rmap_0_address_i                     => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address,                      --             avalon_rmap_slave_0.address
			avs_rmap_0_write_i                       => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write,                        --                                .write
			avs_rmap_0_read_i                        => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read,                         --                                .read
			avs_rmap_0_readdata_o                    => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata,                     --                                .readdata
			avs_rmap_0_writedata_i                   => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata,                    --                                .writedata
			avs_rmap_0_waitrequest_o                 => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest,                  --                                .waitrequest
			rms_rmap_0_wr_address_i                  => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal, --    conduit_end_rmap_mem_slave_0.wr_address_signal
			rms_rmap_0_write_i                       => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,      --                                .write_signal
			rms_rmap_0_writedata_i                   => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,  --                                .writedata_signal
			rms_rmap_0_rd_address_i                  => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal, --                                .rd_address_signal
			rms_rmap_0_read_i                        => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,       --                                .read_signal
			rms_rmap_0_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_0_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_readdata_signal,                       --                                .readdata_signal
			rms_rmap_0_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_0_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_1_wr_address_i                  => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,      --    conduit_end_rmap_mem_slave_1.wr_address_signal
			rms_rmap_1_write_i                       => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,           --                                .write_signal
			rms_rmap_1_writedata_i                   => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,       --                                .writedata_signal
			rms_rmap_1_rd_address_i                  => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,      --                                .rd_address_signal
			rms_rmap_1_read_i                        => communication_module_v2_ch1_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,            --                                .read_signal
			rms_rmap_1_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_1_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_readdata_signal,                       --                                .readdata_signal
			rms_rmap_1_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_1_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_2_wr_address_i                  => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal, --    conduit_end_rmap_mem_slave_2.wr_address_signal
			rms_rmap_2_write_i                       => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,      --                                .write_signal
			rms_rmap_2_writedata_i                   => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,  --                                .writedata_signal
			rms_rmap_2_rd_address_i                  => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal, --                                .rd_address_signal
			rms_rmap_2_read_i                        => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,       --                                .read_signal
			rms_rmap_2_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_2_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_readdata_signal,                       --                                .readdata_signal
			rms_rmap_2_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_2_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_3_wr_address_i                  => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,      --    conduit_end_rmap_mem_slave_3.wr_address_signal
			rms_rmap_3_write_i                       => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,           --                                .write_signal
			rms_rmap_3_writedata_i                   => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,       --                                .writedata_signal
			rms_rmap_3_rd_address_i                  => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,      --                                .rd_address_signal
			rms_rmap_3_read_i                        => communication_module_v2_ch2_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,            --                                .read_signal
			rms_rmap_3_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_3_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_readdata_signal,                       --                                .readdata_signal
			rms_rmap_3_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_3_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_4_wr_address_i                  => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal, --    conduit_end_rmap_mem_slave_4.wr_address_signal
			rms_rmap_4_write_i                       => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,      --                                .write_signal
			rms_rmap_4_writedata_i                   => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,  --                                .writedata_signal
			rms_rmap_4_rd_address_i                  => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal, --                                .rd_address_signal
			rms_rmap_4_read_i                        => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,       --                                .read_signal
			rms_rmap_4_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_4_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_readdata_signal,                       --                                .readdata_signal
			rms_rmap_4_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_4_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_5_wr_address_i                  => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,      --    conduit_end_rmap_mem_slave_5.wr_address_signal
			rms_rmap_5_write_i                       => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,           --                                .write_signal
			rms_rmap_5_writedata_i                   => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,       --                                .writedata_signal
			rms_rmap_5_rd_address_i                  => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,      --                                .rd_address_signal
			rms_rmap_5_read_i                        => communication_module_v2_ch3_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,            --                                .read_signal
			rms_rmap_5_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_5_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_readdata_signal,                       --                                .readdata_signal
			rms_rmap_5_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_5_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_6_wr_address_i                  => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_wr_address_signal, --    conduit_end_rmap_mem_slave_6.wr_address_signal
			rms_rmap_6_write_i                       => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_write_signal,      --                                .write_signal
			rms_rmap_6_writedata_i                   => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_writedata_signal,  --                                .writedata_signal
			rms_rmap_6_rd_address_i                  => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_rd_address_signal, --                                .rd_address_signal
			rms_rmap_6_read_i                        => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_rmap_target_read_signal,       --                                .read_signal
			rms_rmap_6_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_6_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_readdata_signal,                       --                                .readdata_signal
			rms_rmap_6_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_6_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			rms_rmap_7_wr_address_i                  => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_wr_address_signal,      --    conduit_end_rmap_mem_slave_7.wr_address_signal
			rms_rmap_7_write_i                       => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_write_signal,           --                                .write_signal
			rms_rmap_7_writedata_i                   => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_writedata_signal,       --                                .writedata_signal
			rms_rmap_7_rd_address_i                  => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_rd_address_signal,      --                                .rd_address_signal
			rms_rmap_7_read_i                        => communication_module_v2_ch4_conduit_end_rmap_mem_deb_master_fee_hk_read_signal,            --                                .read_signal
			rms_rmap_7_wr_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_wr_waitrequest_signal,                 --                                .wr_waitrequest_signal
			rms_rmap_7_readdata_o                    => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_readdata_signal,                       --                                .readdata_signal
			rms_rmap_7_rd_waitrequest_o              => rmap_mem_ffee_deb_area_conduit_end_rmap_mem_slave_7_rd_waitrequest_signal,                 --                                .rd_waitrequest_signal
			avm_rmap_readdata_i                      => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata,                                     --           avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i                   => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest,                                  --                                .waitrequest
			avm_rmap_address_o                       => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address,                                      --                                .address
			avm_rmap_read_o                          => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read,                                         --                                .read
			avm_rmap_write_o                         => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write,                                        --                                .write
			avm_rmap_writedata_o                     => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata,                                    --                                .writedata
			channel_hk_0_rmap_target_status_i        => communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_status_signal,          --     conduit_end_channel_hk_in_0.rmap_target_status_signal
			channel_hk_0_rmap_target_indicate_i      => communication_module_v2_ch1_conduit_end_channel_hk_out_rmap_target_indicate_signal,        --                                .rmap_target_indicate_signal
			channel_hk_0_spw_link_escape_err_i       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_escape_err_signal,         --                                .spw_link_escape_err_signal
			channel_hk_0_spw_link_credit_err_i       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_credit_err_signal,         --                                .spw_link_credit_err_signal
			channel_hk_0_spw_link_parity_err_i       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_parity_err_signal,         --                                .spw_link_parity_err_signal
			channel_hk_0_spw_link_disconnect_i       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_disconnect_signal,         --                                .spw_link_disconnect_signal
			channel_hk_0_spw_link_started_i          => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_started_signal,            --                                .spw_link_started_signal
			channel_hk_0_spw_link_connecting_i       => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_connecting_signal,         --                                .spw_link_connecting_signal
			channel_hk_0_spw_link_running_i          => communication_module_v2_ch1_conduit_end_channel_hk_out_spw_link_running_signal,            --                                .spw_link_running_signal
			channel_hk_0_frame_counter_i             => communication_module_v2_ch1_conduit_end_channel_hk_out_frame_counter_signal,               --                                .frame_counter_signal
			channel_hk_0_left_buffer_ccd_number_i    => communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,      --                                .left_buffer_ccd_number_signal
			channel_hk_0_right_buffer_ccd_number_i   => communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,     --                                .right_buffer_ccd_number_signal
			channel_hk_0_left_buffer_ccd_side_i      => communication_module_v2_ch1_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,        --                                .left_buffer_ccd_side_signal
			channel_hk_0_right_buffer_ccd_side_i     => communication_module_v2_ch1_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,       --                                .right_buffer_ccd_side_signal
			channel_hk_0_err_left_buffer_overflow_i  => communication_module_v2_ch1_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,    --                                .err_left_buffer_overflow_signal
			channel_hk_0_err_right_buffer_overflow_i => communication_module_v2_ch1_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,   --                                .err_right_buffer_overflow_signal
			channel_hk_1_rmap_target_status_i        => communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_status_signal,          --     conduit_end_channel_hk_in_1.rmap_target_status_signal
			channel_hk_1_rmap_target_indicate_i      => communication_module_v2_ch2_conduit_end_channel_hk_out_rmap_target_indicate_signal,        --                                .rmap_target_indicate_signal
			channel_hk_1_spw_link_escape_err_i       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_escape_err_signal,         --                                .spw_link_escape_err_signal
			channel_hk_1_spw_link_credit_err_i       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_credit_err_signal,         --                                .spw_link_credit_err_signal
			channel_hk_1_spw_link_parity_err_i       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_parity_err_signal,         --                                .spw_link_parity_err_signal
			channel_hk_1_spw_link_disconnect_i       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_disconnect_signal,         --                                .spw_link_disconnect_signal
			channel_hk_1_spw_link_started_i          => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_started_signal,            --                                .spw_link_started_signal
			channel_hk_1_spw_link_connecting_i       => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_connecting_signal,         --                                .spw_link_connecting_signal
			channel_hk_1_spw_link_running_i          => communication_module_v2_ch2_conduit_end_channel_hk_out_spw_link_running_signal,            --                                .spw_link_running_signal
			channel_hk_1_frame_counter_i             => communication_module_v2_ch2_conduit_end_channel_hk_out_frame_counter_signal,               --                                .frame_counter_signal
			channel_hk_1_left_buffer_ccd_number_i    => communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,      --                                .left_buffer_ccd_number_signal
			channel_hk_1_right_buffer_ccd_number_i   => communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,     --                                .right_buffer_ccd_number_signal
			channel_hk_1_left_buffer_ccd_side_i      => communication_module_v2_ch2_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,        --                                .left_buffer_ccd_side_signal
			channel_hk_1_right_buffer_ccd_side_i     => communication_module_v2_ch2_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,       --                                .right_buffer_ccd_side_signal
			channel_hk_1_err_left_buffer_overflow_i  => communication_module_v2_ch2_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,    --                                .err_left_buffer_overflow_signal
			channel_hk_1_err_right_buffer_overflow_i => communication_module_v2_ch2_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,   --                                .err_right_buffer_overflow_signal
			channel_hk_2_rmap_target_status_i        => communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_status_signal,          --     conduit_end_channel_hk_in_2.rmap_target_status_signal
			channel_hk_2_rmap_target_indicate_i      => communication_module_v2_ch3_conduit_end_channel_hk_out_rmap_target_indicate_signal,        --                                .rmap_target_indicate_signal
			channel_hk_2_spw_link_escape_err_i       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_escape_err_signal,         --                                .spw_link_escape_err_signal
			channel_hk_2_spw_link_credit_err_i       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_credit_err_signal,         --                                .spw_link_credit_err_signal
			channel_hk_2_spw_link_parity_err_i       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_parity_err_signal,         --                                .spw_link_parity_err_signal
			channel_hk_2_spw_link_disconnect_i       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_disconnect_signal,         --                                .spw_link_disconnect_signal
			channel_hk_2_spw_link_started_i          => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_started_signal,            --                                .spw_link_started_signal
			channel_hk_2_spw_link_connecting_i       => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_connecting_signal,         --                                .spw_link_connecting_signal
			channel_hk_2_spw_link_running_i          => communication_module_v2_ch3_conduit_end_channel_hk_out_spw_link_running_signal,            --                                .spw_link_running_signal
			channel_hk_2_frame_counter_i             => communication_module_v2_ch3_conduit_end_channel_hk_out_frame_counter_signal,               --                                .frame_counter_signal
			channel_hk_2_left_buffer_ccd_number_i    => communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,      --                                .left_buffer_ccd_number_signal
			channel_hk_2_right_buffer_ccd_number_i   => communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,     --                                .right_buffer_ccd_number_signal
			channel_hk_2_left_buffer_ccd_side_i      => communication_module_v2_ch3_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,        --                                .left_buffer_ccd_side_signal
			channel_hk_2_right_buffer_ccd_side_i     => communication_module_v2_ch3_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,       --                                .right_buffer_ccd_side_signal
			channel_hk_2_err_left_buffer_overflow_i  => communication_module_v2_ch3_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,    --                                .err_left_buffer_overflow_signal
			channel_hk_2_err_right_buffer_overflow_i => communication_module_v2_ch3_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,   --                                .err_right_buffer_overflow_signal
			channel_hk_3_rmap_target_status_i        => communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_status_signal,          --     conduit_end_channel_hk_in_3.rmap_target_status_signal
			channel_hk_3_rmap_target_indicate_i      => communication_module_v2_ch4_conduit_end_channel_hk_out_rmap_target_indicate_signal,        --                                .rmap_target_indicate_signal
			channel_hk_3_spw_link_escape_err_i       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_escape_err_signal,         --                                .spw_link_escape_err_signal
			channel_hk_3_spw_link_credit_err_i       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_credit_err_signal,         --                                .spw_link_credit_err_signal
			channel_hk_3_spw_link_parity_err_i       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_parity_err_signal,         --                                .spw_link_parity_err_signal
			channel_hk_3_spw_link_disconnect_i       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_disconnect_signal,         --                                .spw_link_disconnect_signal
			channel_hk_3_spw_link_started_i          => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_started_signal,            --                                .spw_link_started_signal
			channel_hk_3_spw_link_connecting_i       => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_connecting_signal,         --                                .spw_link_connecting_signal
			channel_hk_3_spw_link_running_i          => communication_module_v2_ch4_conduit_end_channel_hk_out_spw_link_running_signal,            --                                .spw_link_running_signal
			channel_hk_3_frame_counter_i             => communication_module_v2_ch4_conduit_end_channel_hk_out_frame_counter_signal,               --                                .frame_counter_signal
			channel_hk_3_left_buffer_ccd_number_i    => communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_number_signal,      --                                .left_buffer_ccd_number_signal
			channel_hk_3_right_buffer_ccd_number_i   => communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_number_signal,     --                                .right_buffer_ccd_number_signal
			channel_hk_3_left_buffer_ccd_side_i      => communication_module_v2_ch4_conduit_end_channel_hk_out_left_buffer_ccd_side_signal,        --                                .left_buffer_ccd_side_signal
			channel_hk_3_right_buffer_ccd_side_i     => communication_module_v2_ch4_conduit_end_channel_hk_out_right_buffer_ccd_side_signal,       --                                .right_buffer_ccd_side_signal
			channel_hk_3_err_left_buffer_overflow_i  => communication_module_v2_ch4_conduit_end_channel_hk_out_err_left_buffer_overflow_signal,    --                                .err_left_buffer_overflow_signal
			channel_hk_3_err_right_buffer_overflow_i => communication_module_v2_ch4_conduit_end_channel_hk_out_err_right_buffer_overflow_signal,   --                                .err_right_buffer_overflow_signal
			channel_win_mem_addr_offset_i            => communication_module_v2_ch1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal    -- conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
		);

	rs232_uart : component MebX_Qsys_Project_rs232_uart
		port map (
			clk           => clk50_clk,                                       --                 clk.clk
			reset_n       => rst_controller_007_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_2_rs232_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_2_rs232_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_2_rs232_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_2_rs232_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_2_rs232_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_2_rs232_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_2_rs232_uart_s1_readdata,        --                    .readdata
			rxd           => rs232_uart_rxd,                                  -- external_connection.export
			txd           => rs232_uart_txd,                                  --                    .export
			irq           => irq_synchronizer_002_receiver_irq(0)             --                 irq.irq
		);

	rst_controller : component rst_controller_top
		port map (
			clock_sink_clk                          => clk50_clk,                                                                --                  clock_sink.clk
			reset_sink_reset                        => rst_controller_001_reset_out_reset,                                       --                  reset_sink.reset
			reset_source_rs232_reset                => rst_controller_reset_source_rs232_reset,                                  --          reset_source_rs232.reset
			avalon_slave_rst_controller_address     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,     -- avalon_rst_controller_slave.address
			avalon_slave_rst_controller_write       => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,       --                            .write
			avalon_slave_rst_controller_read        => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,        --                            .read
			avalon_slave_rst_controller_writedata   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,   --                            .writedata
			avalon_slave_rst_controller_readdata    => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,    --                            .readdata
			avalon_slave_rst_controller_waitrequest => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest, --                            .waitrequest
			simucam_reset_signal                    => rst_controller_conduit_simucam_reset_t_simucam_reset_signal,              --       conduit_simucam_reset.t_simucam_reset_signal
			reset_input_signal                      => rst_controller_conduit_reset_input_t_reset_input_signal                   --         conduit_reset_input.t_reset_input_signal
		);

	rtcc_alarm : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_rtcc_alarm_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_rtcc_alarm_s1_readdata,     --                    .readdata
			in_port  => rtcc_alarm_export                             -- external_connection.export
		);

	rtcc_cs_n : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_2_rtcc_cs_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_cs_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_cs_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_cs_n_s1_readdata,        --                    .readdata
			out_port   => rtcc_cs_n_export                                -- external_connection.export
		);

	rtcc_sck : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_rtcc_sck_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_sck_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_sck_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_sck_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_sck_s1_readdata,        --                    .readdata
			out_port   => rtcc_sck_export                                -- external_connection.export
		);

	rtcc_sdi : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_rtcc_sdi_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_sdi_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_sdi_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_sdi_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_sdi_s1_readdata,        --                    .readdata
			out_port   => rtcc_sdi_export                                -- external_connection.export
		);

	rtcc_sdo : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_rtcc_sdo_s1_address,        --                  s1.address
			readdata => mm_interconnect_2_rtcc_sdo_s1_readdata,       --                    .readdata
			in_port  => rtcc_sdo_export                               -- external_connection.export
		);

	sd_card_wp_n : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_sd_card_wp_n_s1_address,    --                  s1.address
			readdata => mm_interconnect_2_sd_card_wp_n_s1_readdata,   --                    .readdata
			in_port  => sd_card_wp_n_io_export                        -- external_connection.export
		);

	sync : component sync_ent
		generic map (
			g_SYNC_IRQ_NUMBER     => 11,
			g_PRE_SYNC_IRQ_NUMBER => 12
		)
		port map (
			clock_sink_clk_i                 => clk50_clk,                                          --                     clock.clk
			reset_sink_reset_i               => rst_controller_001_reset_out_reset,                 --                     reset.reset
			avalon_slave_address_i           => mm_interconnect_2_sync_avalon_mm_slave_address,     --           avalon_mm_slave.address
			avalon_slave_read_i              => mm_interconnect_2_sync_avalon_mm_slave_read,        --                          .read
			avalon_slave_write_i             => mm_interconnect_2_sync_avalon_mm_slave_write,       --                          .write
			avalon_slave_writedata_i         => mm_interconnect_2_sync_avalon_mm_slave_writedata,   --                          .writedata
			avalon_slave_readdata_o          => mm_interconnect_2_sync_avalon_mm_slave_readdata,    --                          .readdata
			avalon_slave_waitrequest_o       => mm_interconnect_2_sync_avalon_mm_slave_waitrequest, --                          .waitrequest
			conduit_sync_signal_syncin_en_i  => sync_in_en_conduit,                                 --                sync_in_en.conduit
			conduit_sync_signal_syncout_en_i => sync_out_en_conduit,                                --               sync_out_en.conduit
			conduit_sync_signal_syncin_i     => sync_in_conduit,                                    --                   sync_in.conduit
			conduit_sync_signal_spw1_o       => sync_spw1_conduit,                                  --                 sync_spw1.conduit
			conduit_sync_signal_spw2_o       => sync_spw2_conduit,                                  --                 sync_spw2.conduit
			conduit_sync_signal_spw3_o       => sync_spw3_conduit,                                  --                 sync_spw3.conduit
			conduit_sync_signal_spw4_o       => sync_spw4_conduit,                                  --                 sync_spw4.conduit
			conduit_sync_signal_spw5_o       => sync_spw5_conduit,                                  --                 sync_spw5.conduit
			conduit_sync_signal_spw6_o       => sync_spw6_conduit,                                  --                 sync_spw6.conduit
			conduit_sync_signal_spw7_o       => sync_spw7_conduit,                                  --                 sync_spw7.conduit
			conduit_sync_signal_spw8_o       => sync_spw8_conduit,                                  --                 sync_spw8.conduit
			conduit_sync_signal_syncout_o    => sync_out_conduit,                                   --                  sync_out.conduit
			sync_interrupt_sender_irq_o      => irq_synchronizer_004_receiver_irq(0),               --     sync_interrupt_sender.irq
			pre_sync_interrupt_sender_irq_o  => irq_synchronizer_003_receiver_irq(0)                -- pre_sync_interrupt_sender.irq
		);

	sysid_qsys : component MebX_Qsys_Project_sysid_qsys
		port map (
			clock    => m2_ddr2_memory_afi_half_clk_clk,                       --           clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	temp_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_scl_s1_readdata,        --                    .readdata
			out_port   => temp_scl_export                                -- external_connection.export
		);

	temp_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_sda_s1_readdata,        --                    .readdata
			bidir_port => temp_sda_export                                -- external_connection.export
		);

	timer_1ms : component MebX_Qsys_Project_timer_1ms
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1ms_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1ms_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1ms_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1ms_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1ms_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_receiver_irq(0),               --           irq.irq
			timeout_pulse => timer_1ms_external_port_export                  -- external_port.export
		);

	timer_1us : component MebX_Qsys_Project_timer_1us
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1us_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1us_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1us_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1us_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1us_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_001_receiver_irq(0),           --           irq.irq
			timeout_pulse => timer_1us_external_port_export                  -- external_port.export
		);

	tristate_conduit_bridge_0 : component MebX_Qsys_Project_tristate_conduit_bridge_0
		port map (
			clk                         => m2_ddr2_memory_afi_half_clk_clk,       --   clk.clk
			reset                       => rst_controller_004_reset_out_reset,    -- reset.reset
			request                     => ext_flash_tcm_request,                 --   tcs.request
			grant                       => ext_flash_tcm_grant,                   --      .grant
			tcs_tcm_address_out         => ext_flash_tcm_address_out,             --      .address_out
			tcs_tcm_read_n_out(0)       => ext_flash_tcm_read_n_out,              --      .read_n_out
			tcs_tcm_write_n_out(0)      => ext_flash_tcm_write_n_out,             --      .write_n_out
			tcs_tcm_data_out            => ext_flash_tcm_data_out,                --      .data_out
			tcs_tcm_data_outen          => ext_flash_tcm_data_outen,              --      .data_outen
			tcs_tcm_data_in             => ext_flash_tcm_data_in,                 --      .data_in
			tcs_tcm_chipselect_n_out(0) => ext_flash_tcm_chipselect_n_out,        --      .chipselect_n_out
			tcm_address_out             => tristate_conduit_tcm_address_out,      --   out.tcm_address_out
			tcm_read_n_out              => tristate_conduit_tcm_read_n_out,       --      .tcm_read_n_out
			tcm_write_n_out             => tristate_conduit_tcm_write_n_out,      --      .tcm_write_n_out
			tcm_data_out                => tristate_conduit_tcm_data_out,         --      .tcm_data_out
			tcm_chipselect_n_out        => tristate_conduit_tcm_chipselect_n_out  --      .tcm_chipselect_n_out
		);

	mm_interconnect_0 : component MebX_Qsys_Project_mm_interconnect_0
		port map (
			clk_100_clk_clk                                                       => m2_ddr2_memory_afi_half_clk_clk,                                       --                                               clk_100_clk.clk
			m2_ddr2_memory_afi_clk_clk                                            => m2_ddr2_memory_afi_clk_clk,                                            --                                    m2_ddr2_memory_afi_clk.clk
			m2_ddr2_memory_afi_half_clk_clk                                       => m2_ddr2_memory_afi_half_clk_clk,                                       --                               m2_ddr2_memory_afi_half_clk.clk
			FTDI_UMFT601A_Module_reset_sink_reset_bridge_in_reset_reset           => rst_controller_002_reset_out_reset,                                    --     FTDI_UMFT601A_Module_reset_sink_reset_bridge_in_reset.reset
			m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                                    --            m1_clock_bridge_s0_reset_reset_bridge_in_reset.reset
			m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset       => rst_controller_003_reset_out_reset,                                    -- m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
			m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset                 => rst_controller_003_reset_out_reset,                                    --           m2_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_address      => communication_module_v2_ch1_avalon_mm_left_buffer_master_address,      --  Communication_Module_v2_Ch1_avalon_mm_left_buffer_master.address
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_waitrequest  => communication_module_v2_ch1_avalon_mm_left_buffer_master_waitrequest,  --                                                          .waitrequest
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_read         => communication_module_v2_ch1_avalon_mm_left_buffer_master_read,         --                                                          .read
			Communication_Module_v2_Ch1_avalon_mm_left_buffer_master_readdata     => communication_module_v2_ch1_avalon_mm_left_buffer_master_readdata,     --                                                          .readdata
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_address     => communication_module_v2_ch1_avalon_mm_right_buffer_master_address,     -- Communication_Module_v2_Ch1_avalon_mm_right_buffer_master.address
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_waitrequest => communication_module_v2_ch1_avalon_mm_right_buffer_master_waitrequest, --                                                          .waitrequest
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_read        => communication_module_v2_ch1_avalon_mm_right_buffer_master_read,        --                                                          .read
			Communication_Module_v2_Ch1_avalon_mm_right_buffer_master_readdata    => communication_module_v2_ch1_avalon_mm_right_buffer_master_readdata,    --                                                          .readdata
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_address      => communication_module_v2_ch2_avalon_mm_left_buffer_master_address,      --  Communication_Module_v2_Ch2_avalon_mm_left_buffer_master.address
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_waitrequest  => communication_module_v2_ch2_avalon_mm_left_buffer_master_waitrequest,  --                                                          .waitrequest
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_read         => communication_module_v2_ch2_avalon_mm_left_buffer_master_read,         --                                                          .read
			Communication_Module_v2_Ch2_avalon_mm_left_buffer_master_readdata     => communication_module_v2_ch2_avalon_mm_left_buffer_master_readdata,     --                                                          .readdata
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_address     => communication_module_v2_ch2_avalon_mm_right_buffer_master_address,     -- Communication_Module_v2_Ch2_avalon_mm_right_buffer_master.address
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_waitrequest => communication_module_v2_ch2_avalon_mm_right_buffer_master_waitrequest, --                                                          .waitrequest
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_read        => communication_module_v2_ch2_avalon_mm_right_buffer_master_read,        --                                                          .read
			Communication_Module_v2_Ch2_avalon_mm_right_buffer_master_readdata    => communication_module_v2_ch2_avalon_mm_right_buffer_master_readdata,    --                                                          .readdata
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_address      => communication_module_v2_ch3_avalon_mm_left_buffer_master_address,      --  Communication_Module_v2_Ch3_avalon_mm_left_buffer_master.address
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_waitrequest  => communication_module_v2_ch3_avalon_mm_left_buffer_master_waitrequest,  --                                                          .waitrequest
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_read         => communication_module_v2_ch3_avalon_mm_left_buffer_master_read,         --                                                          .read
			Communication_Module_v2_Ch3_avalon_mm_left_buffer_master_readdata     => communication_module_v2_ch3_avalon_mm_left_buffer_master_readdata,     --                                                          .readdata
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_address     => communication_module_v2_ch3_avalon_mm_right_buffer_master_address,     -- Communication_Module_v2_Ch3_avalon_mm_right_buffer_master.address
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_waitrequest => communication_module_v2_ch3_avalon_mm_right_buffer_master_waitrequest, --                                                          .waitrequest
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_read        => communication_module_v2_ch3_avalon_mm_right_buffer_master_read,        --                                                          .read
			Communication_Module_v2_Ch3_avalon_mm_right_buffer_master_readdata    => communication_module_v2_ch3_avalon_mm_right_buffer_master_readdata,    --                                                          .readdata
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_address      => communication_module_v2_ch4_avalon_mm_left_buffer_master_address,      --  Communication_Module_v2_Ch4_avalon_mm_left_buffer_master.address
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_waitrequest  => communication_module_v2_ch4_avalon_mm_left_buffer_master_waitrequest,  --                                                          .waitrequest
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_read         => communication_module_v2_ch4_avalon_mm_left_buffer_master_read,         --                                                          .read
			Communication_Module_v2_Ch4_avalon_mm_left_buffer_master_readdata     => communication_module_v2_ch4_avalon_mm_left_buffer_master_readdata,     --                                                          .readdata
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_address     => communication_module_v2_ch4_avalon_mm_right_buffer_master_address,     -- Communication_Module_v2_Ch4_avalon_mm_right_buffer_master.address
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_waitrequest => communication_module_v2_ch4_avalon_mm_right_buffer_master_waitrequest, --                                                          .waitrequest
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_read        => communication_module_v2_ch4_avalon_mm_right_buffer_master_read,        --                                                          .read
			Communication_Module_v2_Ch4_avalon_mm_right_buffer_master_readdata    => communication_module_v2_ch4_avalon_mm_right_buffer_master_readdata,    --                                                          .readdata
			ddr2_address_span_extender_expanded_master_address                    => ddr2_address_span_extender_expanded_master_address,                    --                ddr2_address_span_extender_expanded_master.address
			ddr2_address_span_extender_expanded_master_waitrequest                => ddr2_address_span_extender_expanded_master_waitrequest,                --                                                          .waitrequest
			ddr2_address_span_extender_expanded_master_burstcount                 => ddr2_address_span_extender_expanded_master_burstcount,                 --                                                          .burstcount
			ddr2_address_span_extender_expanded_master_byteenable                 => ddr2_address_span_extender_expanded_master_byteenable,                 --                                                          .byteenable
			ddr2_address_span_extender_expanded_master_read                       => ddr2_address_span_extender_expanded_master_read,                       --                                                          .read
			ddr2_address_span_extender_expanded_master_readdata                   => ddr2_address_span_extender_expanded_master_readdata,                   --                                                          .readdata
			ddr2_address_span_extender_expanded_master_readdatavalid              => ddr2_address_span_extender_expanded_master_readdatavalid,              --                                                          .readdatavalid
			ddr2_address_span_extender_expanded_master_write                      => ddr2_address_span_extender_expanded_master_write,                      --                                                          .write
			ddr2_address_span_extender_expanded_master_writedata                  => ddr2_address_span_extender_expanded_master_writedata,                  --                                                          .writedata
			FTDI_UMFT601A_Module_avalon_imgt_master_data_address                  => ftdi_umft601a_module_avalon_imgt_master_data_address,                  --              FTDI_UMFT601A_Module_avalon_imgt_master_data.address
			FTDI_UMFT601A_Module_avalon_imgt_master_data_waitrequest              => ftdi_umft601a_module_avalon_imgt_master_data_waitrequest,              --                                                          .waitrequest
			FTDI_UMFT601A_Module_avalon_imgt_master_data_write                    => ftdi_umft601a_module_avalon_imgt_master_data_write,                    --                                                          .write
			FTDI_UMFT601A_Module_avalon_imgt_master_data_writedata                => ftdi_umft601a_module_avalon_imgt_master_data_writedata,                --                                                          .writedata
			FTDI_UMFT601A_Module_avalon_master_data_address                       => ftdi_umft601a_module_avalon_master_data_address,                       --                   FTDI_UMFT601A_Module_avalon_master_data.address
			FTDI_UMFT601A_Module_avalon_master_data_waitrequest                   => ftdi_umft601a_module_avalon_master_data_waitrequest,                   --                                                          .waitrequest
			FTDI_UMFT601A_Module_avalon_master_data_read                          => ftdi_umft601a_module_avalon_master_data_read,                          --                                                          .read
			FTDI_UMFT601A_Module_avalon_master_data_readdata                      => ftdi_umft601a_module_avalon_master_data_readdata,                      --                                                          .readdata
			FTDI_UMFT601A_Module_avalon_master_data_write                         => ftdi_umft601a_module_avalon_master_data_write,                         --                                                          .write
			FTDI_UMFT601A_Module_avalon_master_data_writedata                     => ftdi_umft601a_module_avalon_master_data_writedata,                     --                                                          .writedata
			Memory_Filler_avalon_master_data_address                              => memory_filler_avalon_master_data_address,                              --                          Memory_Filler_avalon_master_data.address
			Memory_Filler_avalon_master_data_waitrequest                          => memory_filler_avalon_master_data_waitrequest,                          --                                                          .waitrequest
			Memory_Filler_avalon_master_data_write                                => memory_filler_avalon_master_data_write,                                --                                                          .write
			Memory_Filler_avalon_master_data_writedata                            => memory_filler_avalon_master_data_writedata,                            --                                                          .writedata
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address                  => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_address,                  --              rmap_mem_ffee_deb_area_avalon_mm_rmap_master.address
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest              => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_waitrequest,              --                                                          .waitrequest
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read                     => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_read,                     --                                                          .read
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata                 => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_readdata,                 --                                                          .readdata
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write                    => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_write,                    --                                                          .write
			rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata                => rmap_mem_ffee_deb_area_avalon_mm_rmap_master_writedata,                --                                                          .writedata
			m1_clock_bridge_s0_address                                            => mm_interconnect_0_m1_clock_bridge_s0_address,                          --                                        m1_clock_bridge_s0.address
			m1_clock_bridge_s0_write                                              => mm_interconnect_0_m1_clock_bridge_s0_write,                            --                                                          .write
			m1_clock_bridge_s0_read                                               => mm_interconnect_0_m1_clock_bridge_s0_read,                             --                                                          .read
			m1_clock_bridge_s0_readdata                                           => mm_interconnect_0_m1_clock_bridge_s0_readdata,                         --                                                          .readdata
			m1_clock_bridge_s0_writedata                                          => mm_interconnect_0_m1_clock_bridge_s0_writedata,                        --                                                          .writedata
			m1_clock_bridge_s0_burstcount                                         => mm_interconnect_0_m1_clock_bridge_s0_burstcount,                       --                                                          .burstcount
			m1_clock_bridge_s0_byteenable                                         => mm_interconnect_0_m1_clock_bridge_s0_byteenable,                       --                                                          .byteenable
			m1_clock_bridge_s0_readdatavalid                                      => mm_interconnect_0_m1_clock_bridge_s0_readdatavalid,                    --                                                          .readdatavalid
			m1_clock_bridge_s0_waitrequest                                        => mm_interconnect_0_m1_clock_bridge_s0_waitrequest,                      --                                                          .waitrequest
			m1_clock_bridge_s0_debugaccess                                        => mm_interconnect_0_m1_clock_bridge_s0_debugaccess,                      --                                                          .debugaccess
			m2_ddr2_memory_avl_address                                            => mm_interconnect_0_m2_ddr2_memory_avl_address,                          --                                        m2_ddr2_memory_avl.address
			m2_ddr2_memory_avl_write                                              => mm_interconnect_0_m2_ddr2_memory_avl_write,                            --                                                          .write
			m2_ddr2_memory_avl_read                                               => mm_interconnect_0_m2_ddr2_memory_avl_read,                             --                                                          .read
			m2_ddr2_memory_avl_readdata                                           => mm_interconnect_0_m2_ddr2_memory_avl_readdata,                         --                                                          .readdata
			m2_ddr2_memory_avl_writedata                                          => mm_interconnect_0_m2_ddr2_memory_avl_writedata,                        --                                                          .writedata
			m2_ddr2_memory_avl_beginbursttransfer                                 => mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer,               --                                                          .beginbursttransfer
			m2_ddr2_memory_avl_burstcount                                         => mm_interconnect_0_m2_ddr2_memory_avl_burstcount,                       --                                                          .burstcount
			m2_ddr2_memory_avl_byteenable                                         => mm_interconnect_0_m2_ddr2_memory_avl_byteenable,                       --                                                          .byteenable
			m2_ddr2_memory_avl_readdatavalid                                      => mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid,                    --                                                          .readdatavalid
			m2_ddr2_memory_avl_waitrequest                                        => mm_interconnect_0_m2_ddr2_memory_avl_inv                               --                                                          .waitrequest
		);

	mm_interconnect_1 : component MebX_Qsys_Project_mm_interconnect_1
		port map (
			clk_100_clk_clk                                                => m2_ddr2_memory_afi_half_clk_clk,                                                  --                                        clk_100_clk.clk
			ext_flash_reset_reset_bridge_in_reset_reset                    => rst_controller_004_reset_out_reset,                                               --              ext_flash_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                                               --            jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                 => rst_controller_006_reset_out_reset,                                               --           nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                               => nios2_gen2_0_data_master_address,                                                 --                           nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                           => nios2_gen2_0_data_master_waitrequest,                                             --                                                   .waitrequest
			nios2_gen2_0_data_master_byteenable                            => nios2_gen2_0_data_master_byteenable,                                              --                                                   .byteenable
			nios2_gen2_0_data_master_read                                  => nios2_gen2_0_data_master_read,                                                    --                                                   .read
			nios2_gen2_0_data_master_readdata                              => nios2_gen2_0_data_master_readdata,                                                --                                                   .readdata
			nios2_gen2_0_data_master_write                                 => nios2_gen2_0_data_master_write,                                                   --                                                   .write
			nios2_gen2_0_data_master_writedata                             => nios2_gen2_0_data_master_writedata,                                               --                                                   .writedata
			nios2_gen2_0_data_master_debugaccess                           => nios2_gen2_0_data_master_debugaccess,                                             --                                                   .debugaccess
			nios2_gen2_0_instruction_master_address                        => nios2_gen2_0_instruction_master_address,                                          --                    nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                    => nios2_gen2_0_instruction_master_waitrequest,                                      --                                                   .waitrequest
			nios2_gen2_0_instruction_master_burstcount                     => nios2_gen2_0_instruction_master_burstcount,                                       --                                                   .burstcount
			nios2_gen2_0_instruction_master_read                           => nios2_gen2_0_instruction_master_read,                                             --                                                   .read
			nios2_gen2_0_instruction_master_readdata                       => nios2_gen2_0_instruction_master_readdata,                                         --                                                   .readdata
			nios2_gen2_0_instruction_master_readdatavalid                  => nios2_gen2_0_instruction_master_readdatavalid,                                    --                                                   .readdatavalid
			clock_bridge_afi_50_s0_address                                 => mm_interconnect_1_clock_bridge_afi_50_s0_address,                                 --                             clock_bridge_afi_50_s0.address
			clock_bridge_afi_50_s0_write                                   => mm_interconnect_1_clock_bridge_afi_50_s0_write,                                   --                                                   .write
			clock_bridge_afi_50_s0_read                                    => mm_interconnect_1_clock_bridge_afi_50_s0_read,                                    --                                                   .read
			clock_bridge_afi_50_s0_readdata                                => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,                                --                                                   .readdata
			clock_bridge_afi_50_s0_writedata                               => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,                               --                                                   .writedata
			clock_bridge_afi_50_s0_burstcount                              => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,                              --                                                   .burstcount
			clock_bridge_afi_50_s0_byteenable                              => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,                              --                                                   .byteenable
			clock_bridge_afi_50_s0_readdatavalid                           => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid,                           --                                                   .readdatavalid
			clock_bridge_afi_50_s0_waitrequest                             => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,                             --                                                   .waitrequest
			clock_bridge_afi_50_s0_debugaccess                             => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,                             --                                                   .debugaccess
			Communication_Module_v2_Ch1_avalon_mm_config_slave_address     => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_address,     -- Communication_Module_v2_Ch1_avalon_mm_config_slave.address
			Communication_Module_v2_Ch1_avalon_mm_config_slave_write       => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_write,       --                                                   .write
			Communication_Module_v2_Ch1_avalon_mm_config_slave_read        => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_read,        --                                                   .read
			Communication_Module_v2_Ch1_avalon_mm_config_slave_readdata    => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_readdata,    --                                                   .readdata
			Communication_Module_v2_Ch1_avalon_mm_config_slave_writedata   => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_writedata,   --                                                   .writedata
			Communication_Module_v2_Ch1_avalon_mm_config_slave_waitrequest => mm_interconnect_1_communication_module_v2_ch1_avalon_mm_config_slave_waitrequest, --                                                   .waitrequest
			Communication_Module_v2_Ch2_avalon_mm_config_slave_address     => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_address,     -- Communication_Module_v2_Ch2_avalon_mm_config_slave.address
			Communication_Module_v2_Ch2_avalon_mm_config_slave_write       => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_write,       --                                                   .write
			Communication_Module_v2_Ch2_avalon_mm_config_slave_read        => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_read,        --                                                   .read
			Communication_Module_v2_Ch2_avalon_mm_config_slave_readdata    => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_readdata,    --                                                   .readdata
			Communication_Module_v2_Ch2_avalon_mm_config_slave_writedata   => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_writedata,   --                                                   .writedata
			Communication_Module_v2_Ch2_avalon_mm_config_slave_waitrequest => mm_interconnect_1_communication_module_v2_ch2_avalon_mm_config_slave_waitrequest, --                                                   .waitrequest
			Communication_Module_v2_Ch3_avalon_mm_config_slave_address     => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_address,     -- Communication_Module_v2_Ch3_avalon_mm_config_slave.address
			Communication_Module_v2_Ch3_avalon_mm_config_slave_write       => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_write,       --                                                   .write
			Communication_Module_v2_Ch3_avalon_mm_config_slave_read        => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_read,        --                                                   .read
			Communication_Module_v2_Ch3_avalon_mm_config_slave_readdata    => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_readdata,    --                                                   .readdata
			Communication_Module_v2_Ch3_avalon_mm_config_slave_writedata   => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_writedata,   --                                                   .writedata
			Communication_Module_v2_Ch3_avalon_mm_config_slave_waitrequest => mm_interconnect_1_communication_module_v2_ch3_avalon_mm_config_slave_waitrequest, --                                                   .waitrequest
			Communication_Module_v2_Ch4_avalon_mm_config_slave_address     => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_address,     -- Communication_Module_v2_Ch4_avalon_mm_config_slave.address
			Communication_Module_v2_Ch4_avalon_mm_config_slave_write       => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_write,       --                                                   .write
			Communication_Module_v2_Ch4_avalon_mm_config_slave_read        => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_read,        --                                                   .read
			Communication_Module_v2_Ch4_avalon_mm_config_slave_readdata    => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_readdata,    --                                                   .readdata
			Communication_Module_v2_Ch4_avalon_mm_config_slave_writedata   => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_writedata,   --                                                   .writedata
			Communication_Module_v2_Ch4_avalon_mm_config_slave_waitrequest => mm_interconnect_1_communication_module_v2_ch4_avalon_mm_config_slave_waitrequest, --                                                   .waitrequest
			ddr2_address_span_extender_cntl_write                          => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                          --                    ddr2_address_span_extender_cntl.write
			ddr2_address_span_extender_cntl_read                           => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                           --                                                   .read
			ddr2_address_span_extender_cntl_readdata                       => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                       --                                                   .readdata
			ddr2_address_span_extender_cntl_writedata                      => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,                      --                                                   .writedata
			ddr2_address_span_extender_cntl_byteenable                     => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,                     --                                                   .byteenable
			ddr2_address_span_extender_windowed_slave_address              => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,              --          ddr2_address_span_extender_windowed_slave.address
			ddr2_address_span_extender_windowed_slave_write                => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,                --                                                   .write
			ddr2_address_span_extender_windowed_slave_read                 => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,                 --                                                   .read
			ddr2_address_span_extender_windowed_slave_readdata             => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,             --                                                   .readdata
			ddr2_address_span_extender_windowed_slave_writedata            => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,            --                                                   .writedata
			ddr2_address_span_extender_windowed_slave_burstcount           => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,           --                                                   .burstcount
			ddr2_address_span_extender_windowed_slave_byteenable           => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,           --                                                   .byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid        => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid,        --                                                   .readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,          --                                                   .waitrequest
			ext_flash_uas_address                                          => mm_interconnect_1_ext_flash_uas_address,                                          --                                      ext_flash_uas.address
			ext_flash_uas_write                                            => mm_interconnect_1_ext_flash_uas_write,                                            --                                                   .write
			ext_flash_uas_read                                             => mm_interconnect_1_ext_flash_uas_read,                                             --                                                   .read
			ext_flash_uas_readdata                                         => mm_interconnect_1_ext_flash_uas_readdata,                                         --                                                   .readdata
			ext_flash_uas_writedata                                        => mm_interconnect_1_ext_flash_uas_writedata,                                        --                                                   .writedata
			ext_flash_uas_burstcount                                       => mm_interconnect_1_ext_flash_uas_burstcount,                                       --                                                   .burstcount
			ext_flash_uas_byteenable                                       => mm_interconnect_1_ext_flash_uas_byteenable,                                       --                                                   .byteenable
			ext_flash_uas_readdatavalid                                    => mm_interconnect_1_ext_flash_uas_readdatavalid,                                    --                                                   .readdatavalid
			ext_flash_uas_waitrequest                                      => mm_interconnect_1_ext_flash_uas_waitrequest,                                      --                                                   .waitrequest
			ext_flash_uas_lock                                             => mm_interconnect_1_ext_flash_uas_lock,                                             --                                                   .lock
			ext_flash_uas_debugaccess                                      => mm_interconnect_1_ext_flash_uas_debugaccess,                                      --                                                   .debugaccess
			FTDI_UMFT601A_Module_avalon_slave_config_address               => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_address,               --           FTDI_UMFT601A_Module_avalon_slave_config.address
			FTDI_UMFT601A_Module_avalon_slave_config_write                 => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_write,                 --                                                   .write
			FTDI_UMFT601A_Module_avalon_slave_config_read                  => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_read,                  --                                                   .read
			FTDI_UMFT601A_Module_avalon_slave_config_readdata              => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_readdata,              --                                                   .readdata
			FTDI_UMFT601A_Module_avalon_slave_config_writedata             => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_writedata,             --                                                   .writedata
			FTDI_UMFT601A_Module_avalon_slave_config_waitrequest           => mm_interconnect_1_ftdi_umft601a_module_avalon_slave_config_waitrequest,           --                                                   .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                          => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address,                          --                      jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                            => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write,                            --                                                   .write
			jtag_uart_0_avalon_jtag_slave_read                             => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read,                             --                                                   .read
			jtag_uart_0_avalon_jtag_slave_readdata                         => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,                         --                                                   .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                        => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,                        --                                                   .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,                      --                                                   .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                       => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,                       --                                                   .chipselect
			Memory_Filler_avalon_slave_config_address                      => mm_interconnect_1_memory_filler_avalon_slave_config_address,                      --                  Memory_Filler_avalon_slave_config.address
			Memory_Filler_avalon_slave_config_write                        => mm_interconnect_1_memory_filler_avalon_slave_config_write,                        --                                                   .write
			Memory_Filler_avalon_slave_config_read                         => mm_interconnect_1_memory_filler_avalon_slave_config_read,                         --                                                   .read
			Memory_Filler_avalon_slave_config_readdata                     => mm_interconnect_1_memory_filler_avalon_slave_config_readdata,                     --                                                   .readdata
			Memory_Filler_avalon_slave_config_writedata                    => mm_interconnect_1_memory_filler_avalon_slave_config_writedata,                    --                                                   .writedata
			Memory_Filler_avalon_slave_config_byteenable                   => mm_interconnect_1_memory_filler_avalon_slave_config_byteenable,                   --                                                   .byteenable
			Memory_Filler_avalon_slave_config_waitrequest                  => mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest,                  --                                                   .waitrequest
			nios2_gen2_0_debug_mem_slave_address                           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,                           --                       nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,                             --                                                   .write
			nios2_gen2_0_debug_mem_slave_read                              => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,                              --                                                   .read
			nios2_gen2_0_debug_mem_slave_readdata                          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,                          --                                                   .readdata
			nios2_gen2_0_debug_mem_slave_writedata                         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,                         --                                                   .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                        => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,                        --                                                   .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest,                       --                                                   .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess,                       --                                                   .debugaccess
			onchip_memory_s1_address                                       => mm_interconnect_1_onchip_memory_s1_address,                                       --                                   onchip_memory_s1.address
			onchip_memory_s1_write                                         => mm_interconnect_1_onchip_memory_s1_write,                                         --                                                   .write
			onchip_memory_s1_readdata                                      => mm_interconnect_1_onchip_memory_s1_readdata,                                      --                                                   .readdata
			onchip_memory_s1_writedata                                     => mm_interconnect_1_onchip_memory_s1_writedata,                                     --                                                   .writedata
			onchip_memory_s1_byteenable                                    => mm_interconnect_1_onchip_memory_s1_byteenable,                                    --                                                   .byteenable
			onchip_memory_s1_chipselect                                    => mm_interconnect_1_onchip_memory_s1_chipselect,                                    --                                                   .chipselect
			onchip_memory_s1_clken                                         => mm_interconnect_1_onchip_memory_s1_clken,                                         --                                                   .clken
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address           => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_address,           --       rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0.address
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write             => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_write,             --                                                   .write
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read              => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_read,              --                                                   .read
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata          => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_readdata,          --                                                   .readdata
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata         => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_writedata,         --                                                   .writedata
			rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest       => mm_interconnect_1_rmap_mem_ffee_aeb_1_area_avalon_rmap_slave_0_waitrequest,       --                                                   .waitrequest
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address           => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_address,           --       rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0.address
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write             => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_write,             --                                                   .write
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read              => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_read,              --                                                   .read
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata          => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_readdata,          --                                                   .readdata
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata         => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_writedata,         --                                                   .writedata
			rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest       => mm_interconnect_1_rmap_mem_ffee_aeb_2_area_avalon_rmap_slave_0_waitrequest,       --                                                   .waitrequest
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address           => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_address,           --       rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0.address
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write             => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_write,             --                                                   .write
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read              => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_read,              --                                                   .read
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata          => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_readdata,          --                                                   .readdata
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata         => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_writedata,         --                                                   .writedata
			rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest       => mm_interconnect_1_rmap_mem_ffee_aeb_3_area_avalon_rmap_slave_0_waitrequest,       --                                                   .waitrequest
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address           => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_address,           --       rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0.address
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write             => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_write,             --                                                   .write
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read              => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_read,              --                                                   .read
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata          => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_readdata,          --                                                   .readdata
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata         => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_writedata,         --                                                   .writedata
			rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest       => mm_interconnect_1_rmap_mem_ffee_aeb_4_area_avalon_rmap_slave_0_waitrequest,       --                                                   .waitrequest
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address             => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_address,             --         rmap_mem_ffee_deb_area_avalon_rmap_slave_0.address
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write               => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_write,               --                                                   .write
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read                => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_read,                --                                                   .read
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata            => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_readdata,            --                                                   .readdata
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata           => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_writedata,           --                                                   .writedata
			rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest         => mm_interconnect_1_rmap_mem_ffee_deb_area_avalon_rmap_slave_0_waitrequest,         --                                                   .waitrequest
			sysid_qsys_control_slave_address                               => mm_interconnect_1_sysid_qsys_control_slave_address,                               --                           sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                              => mm_interconnect_1_sysid_qsys_control_slave_readdata                               --                                                   .readdata
		);

	mm_interconnect_2 : component MebX_Qsys_Project_mm_interconnect_2
		port map (
			clk_50_clk_clk                                                       => clk50_clk,                                                                              --                                               clk_50_clk.clk
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset             => rst_controller_001_reset_out_reset,                                                     --       clock_bridge_afi_50_m0_reset_reset_bridge_in_reset.reset
			rs232_uart_reset_reset_bridge_in_reset_reset                         => rst_controller_007_reset_out_reset,                                                     --                   rs232_uart_reset_reset_bridge_in_reset.reset
			clock_bridge_afi_50_m0_address                                       => clock_bridge_afi_50_m0_address,                                                         --                                   clock_bridge_afi_50_m0.address
			clock_bridge_afi_50_m0_waitrequest                                   => clock_bridge_afi_50_m0_waitrequest,                                                     --                                                         .waitrequest
			clock_bridge_afi_50_m0_burstcount                                    => clock_bridge_afi_50_m0_burstcount,                                                      --                                                         .burstcount
			clock_bridge_afi_50_m0_byteenable                                    => clock_bridge_afi_50_m0_byteenable,                                                      --                                                         .byteenable
			clock_bridge_afi_50_m0_read                                          => clock_bridge_afi_50_m0_read,                                                            --                                                         .read
			clock_bridge_afi_50_m0_readdata                                      => clock_bridge_afi_50_m0_readdata,                                                        --                                                         .readdata
			clock_bridge_afi_50_m0_readdatavalid                                 => clock_bridge_afi_50_m0_readdatavalid,                                                   --                                                         .readdatavalid
			clock_bridge_afi_50_m0_write                                         => clock_bridge_afi_50_m0_write,                                                           --                                                         .write
			clock_bridge_afi_50_m0_writedata                                     => clock_bridge_afi_50_m0_writedata,                                                       --                                                         .writedata
			clock_bridge_afi_50_m0_debugaccess                                   => clock_bridge_afi_50_m0_debugaccess,                                                     --                                                         .debugaccess
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                                                         .write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                                                         .read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                                                         .readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                                                         .writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                                                         .byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                                                         .waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  --                                                         .chipselect
			csense_adc_fo_s1_address                                             => mm_interconnect_2_csense_adc_fo_s1_address,                                             --                                         csense_adc_fo_s1.address
			csense_adc_fo_s1_write                                               => mm_interconnect_2_csense_adc_fo_s1_write,                                               --                                                         .write
			csense_adc_fo_s1_readdata                                            => mm_interconnect_2_csense_adc_fo_s1_readdata,                                            --                                                         .readdata
			csense_adc_fo_s1_writedata                                           => mm_interconnect_2_csense_adc_fo_s1_writedata,                                           --                                                         .writedata
			csense_adc_fo_s1_chipselect                                          => mm_interconnect_2_csense_adc_fo_s1_chipselect,                                          --                                                         .chipselect
			csense_cs_n_s1_address                                               => mm_interconnect_2_csense_cs_n_s1_address,                                               --                                           csense_cs_n_s1.address
			csense_cs_n_s1_write                                                 => mm_interconnect_2_csense_cs_n_s1_write,                                                 --                                                         .write
			csense_cs_n_s1_readdata                                              => mm_interconnect_2_csense_cs_n_s1_readdata,                                              --                                                         .readdata
			csense_cs_n_s1_writedata                                             => mm_interconnect_2_csense_cs_n_s1_writedata,                                             --                                                         .writedata
			csense_cs_n_s1_chipselect                                            => mm_interconnect_2_csense_cs_n_s1_chipselect,                                            --                                                         .chipselect
			csense_sck_s1_address                                                => mm_interconnect_2_csense_sck_s1_address,                                                --                                            csense_sck_s1.address
			csense_sck_s1_write                                                  => mm_interconnect_2_csense_sck_s1_write,                                                  --                                                         .write
			csense_sck_s1_readdata                                               => mm_interconnect_2_csense_sck_s1_readdata,                                               --                                                         .readdata
			csense_sck_s1_writedata                                              => mm_interconnect_2_csense_sck_s1_writedata,                                              --                                                         .writedata
			csense_sck_s1_chipselect                                             => mm_interconnect_2_csense_sck_s1_chipselect,                                             --                                                         .chipselect
			csense_sdi_s1_address                                                => mm_interconnect_2_csense_sdi_s1_address,                                                --                                            csense_sdi_s1.address
			csense_sdi_s1_write                                                  => mm_interconnect_2_csense_sdi_s1_write,                                                  --                                                         .write
			csense_sdi_s1_readdata                                               => mm_interconnect_2_csense_sdi_s1_readdata,                                               --                                                         .readdata
			csense_sdi_s1_writedata                                              => mm_interconnect_2_csense_sdi_s1_writedata,                                              --                                                         .writedata
			csense_sdi_s1_chipselect                                             => mm_interconnect_2_csense_sdi_s1_chipselect,                                             --                                                         .chipselect
			csense_sdo_s1_address                                                => mm_interconnect_2_csense_sdo_s1_address,                                                --                                            csense_sdo_s1.address
			csense_sdo_s1_readdata                                               => mm_interconnect_2_csense_sdo_s1_readdata,                                               --                                                         .readdata
			m1_ddr2_i2c_scl_s1_address                                           => mm_interconnect_2_m1_ddr2_i2c_scl_s1_address,                                           --                                       m1_ddr2_i2c_scl_s1.address
			m1_ddr2_i2c_scl_s1_write                                             => mm_interconnect_2_m1_ddr2_i2c_scl_s1_write,                                             --                                                         .write
			m1_ddr2_i2c_scl_s1_readdata                                          => mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata,                                          --                                                         .readdata
			m1_ddr2_i2c_scl_s1_writedata                                         => mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata,                                         --                                                         .writedata
			m1_ddr2_i2c_scl_s1_chipselect                                        => mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect,                                        --                                                         .chipselect
			m1_ddr2_i2c_sda_s1_address                                           => mm_interconnect_2_m1_ddr2_i2c_sda_s1_address,                                           --                                       m1_ddr2_i2c_sda_s1.address
			m1_ddr2_i2c_sda_s1_write                                             => mm_interconnect_2_m1_ddr2_i2c_sda_s1_write,                                             --                                                         .write
			m1_ddr2_i2c_sda_s1_readdata                                          => mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata,                                          --                                                         .readdata
			m1_ddr2_i2c_sda_s1_writedata                                         => mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata,                                         --                                                         .writedata
			m1_ddr2_i2c_sda_s1_chipselect                                        => mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect,                                        --                                                         .chipselect
			m2_ddr2_i2c_scl_s1_address                                           => mm_interconnect_2_m2_ddr2_i2c_scl_s1_address,                                           --                                       m2_ddr2_i2c_scl_s1.address
			m2_ddr2_i2c_scl_s1_write                                             => mm_interconnect_2_m2_ddr2_i2c_scl_s1_write,                                             --                                                         .write
			m2_ddr2_i2c_scl_s1_readdata                                          => mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata,                                          --                                                         .readdata
			m2_ddr2_i2c_scl_s1_writedata                                         => mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata,                                         --                                                         .writedata
			m2_ddr2_i2c_scl_s1_chipselect                                        => mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect,                                        --                                                         .chipselect
			m2_ddr2_i2c_sda_s1_address                                           => mm_interconnect_2_m2_ddr2_i2c_sda_s1_address,                                           --                                       m2_ddr2_i2c_sda_s1.address
			m2_ddr2_i2c_sda_s1_write                                             => mm_interconnect_2_m2_ddr2_i2c_sda_s1_write,                                             --                                                         .write
			m2_ddr2_i2c_sda_s1_readdata                                          => mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata,                                          --                                                         .readdata
			m2_ddr2_i2c_sda_s1_writedata                                         => mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata,                                         --                                                         .writedata
			m2_ddr2_i2c_sda_s1_chipselect                                        => mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect,                                        --                                                         .chipselect
			pio_BUTTON_s1_address                                                => mm_interconnect_2_pio_button_s1_address,                                                --                                            pio_BUTTON_s1.address
			pio_BUTTON_s1_readdata                                               => mm_interconnect_2_pio_button_s1_readdata,                                               --                                                         .readdata
			pio_ctrl_io_lvds_s1_address                                          => mm_interconnect_2_pio_ctrl_io_lvds_s1_address,                                          --                                      pio_ctrl_io_lvds_s1.address
			pio_ctrl_io_lvds_s1_write                                            => mm_interconnect_2_pio_ctrl_io_lvds_s1_write,                                            --                                                         .write
			pio_ctrl_io_lvds_s1_readdata                                         => mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata,                                         --                                                         .readdata
			pio_ctrl_io_lvds_s1_writedata                                        => mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata,                                        --                                                         .writedata
			pio_ctrl_io_lvds_s1_chipselect                                       => mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect,                                       --                                                         .chipselect
			pio_DIP_s1_address                                                   => mm_interconnect_2_pio_dip_s1_address,                                                   --                                               pio_DIP_s1.address
			pio_DIP_s1_readdata                                                  => mm_interconnect_2_pio_dip_s1_readdata,                                                  --                                                         .readdata
			pio_EXT_s1_address                                                   => mm_interconnect_2_pio_ext_s1_address,                                                   --                                               pio_EXT_s1.address
			pio_EXT_s1_readdata                                                  => mm_interconnect_2_pio_ext_s1_readdata,                                                  --                                                         .readdata
			pio_ftdi_umft601a_module_reset_s1_address                            => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_address,                            --                        pio_ftdi_umft601a_module_reset_s1.address
			pio_ftdi_umft601a_module_reset_s1_write                              => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write,                              --                                                         .write
			pio_ftdi_umft601a_module_reset_s1_readdata                           => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_readdata,                           --                                                         .readdata
			pio_ftdi_umft601a_module_reset_s1_writedata                          => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_writedata,                          --                                                         .writedata
			pio_ftdi_umft601a_module_reset_s1_chipselect                         => mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_chipselect,                         --                                                         .chipselect
			pio_iso_logic_signal_enable_s1_address                               => mm_interconnect_2_pio_iso_logic_signal_enable_s1_address,                               --                           pio_iso_logic_signal_enable_s1.address
			pio_iso_logic_signal_enable_s1_write                                 => mm_interconnect_2_pio_iso_logic_signal_enable_s1_write,                                 --                                                         .write
			pio_iso_logic_signal_enable_s1_readdata                              => mm_interconnect_2_pio_iso_logic_signal_enable_s1_readdata,                              --                                                         .readdata
			pio_iso_logic_signal_enable_s1_writedata                             => mm_interconnect_2_pio_iso_logic_signal_enable_s1_writedata,                             --                                                         .writedata
			pio_iso_logic_signal_enable_s1_chipselect                            => mm_interconnect_2_pio_iso_logic_signal_enable_s1_chipselect,                            --                                                         .chipselect
			pio_LED_s1_address                                                   => mm_interconnect_2_pio_led_s1_address,                                                   --                                               pio_LED_s1.address
			pio_LED_s1_write                                                     => mm_interconnect_2_pio_led_s1_write,                                                     --                                                         .write
			pio_LED_s1_readdata                                                  => mm_interconnect_2_pio_led_s1_readdata,                                                  --                                                         .readdata
			pio_LED_s1_writedata                                                 => mm_interconnect_2_pio_led_s1_writedata,                                                 --                                                         .writedata
			pio_LED_s1_chipselect                                                => mm_interconnect_2_pio_led_s1_chipselect,                                                --                                                         .chipselect
			pio_LED_painel_s1_address                                            => mm_interconnect_2_pio_led_painel_s1_address,                                            --                                        pio_LED_painel_s1.address
			pio_LED_painel_s1_write                                              => mm_interconnect_2_pio_led_painel_s1_write,                                              --                                                         .write
			pio_LED_painel_s1_readdata                                           => mm_interconnect_2_pio_led_painel_s1_readdata,                                           --                                                         .readdata
			pio_LED_painel_s1_writedata                                          => mm_interconnect_2_pio_led_painel_s1_writedata,                                          --                                                         .writedata
			pio_LED_painel_s1_chipselect                                         => mm_interconnect_2_pio_led_painel_s1_chipselect,                                         --                                                         .chipselect
			pio_spw_demux_ch_1_select_s1_address                                 => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_address,                                 --                             pio_spw_demux_ch_1_select_s1.address
			pio_spw_demux_ch_1_select_s1_write                                   => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write,                                   --                                                         .write
			pio_spw_demux_ch_1_select_s1_readdata                                => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_readdata,                                --                                                         .readdata
			pio_spw_demux_ch_1_select_s1_writedata                               => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_writedata,                               --                                                         .writedata
			pio_spw_demux_ch_1_select_s1_chipselect                              => mm_interconnect_2_pio_spw_demux_ch_1_select_s1_chipselect,                              --                                                         .chipselect
			pio_spw_demux_ch_2_select_s1_address                                 => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_address,                                 --                             pio_spw_demux_ch_2_select_s1.address
			pio_spw_demux_ch_2_select_s1_write                                   => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write,                                   --                                                         .write
			pio_spw_demux_ch_2_select_s1_readdata                                => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_readdata,                                --                                                         .readdata
			pio_spw_demux_ch_2_select_s1_writedata                               => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_writedata,                               --                                                         .writedata
			pio_spw_demux_ch_2_select_s1_chipselect                              => mm_interconnect_2_pio_spw_demux_ch_2_select_s1_chipselect,                              --                                                         .chipselect
			pio_spw_demux_ch_3_select_s1_address                                 => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_address,                                 --                             pio_spw_demux_ch_3_select_s1.address
			pio_spw_demux_ch_3_select_s1_write                                   => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write,                                   --                                                         .write
			pio_spw_demux_ch_3_select_s1_readdata                                => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_readdata,                                --                                                         .readdata
			pio_spw_demux_ch_3_select_s1_writedata                               => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_writedata,                               --                                                         .writedata
			pio_spw_demux_ch_3_select_s1_chipselect                              => mm_interconnect_2_pio_spw_demux_ch_3_select_s1_chipselect,                              --                                                         .chipselect
			pio_spw_demux_ch_4_select_s1_address                                 => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_address,                                 --                             pio_spw_demux_ch_4_select_s1.address
			pio_spw_demux_ch_4_select_s1_write                                   => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write,                                   --                                                         .write
			pio_spw_demux_ch_4_select_s1_readdata                                => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_readdata,                                --                                                         .readdata
			pio_spw_demux_ch_4_select_s1_writedata                               => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_writedata,                               --                                                         .writedata
			pio_spw_demux_ch_4_select_s1_chipselect                              => mm_interconnect_2_pio_spw_demux_ch_4_select_s1_chipselect,                              --                                                         .chipselect
			rs232_uart_s1_address                                                => mm_interconnect_2_rs232_uart_s1_address,                                                --                                            rs232_uart_s1.address
			rs232_uart_s1_write                                                  => mm_interconnect_2_rs232_uart_s1_write,                                                  --                                                         .write
			rs232_uart_s1_read                                                   => mm_interconnect_2_rs232_uart_s1_read,                                                   --                                                         .read
			rs232_uart_s1_readdata                                               => mm_interconnect_2_rs232_uart_s1_readdata,                                               --                                                         .readdata
			rs232_uart_s1_writedata                                              => mm_interconnect_2_rs232_uart_s1_writedata,                                              --                                                         .writedata
			rs232_uart_s1_begintransfer                                          => mm_interconnect_2_rs232_uart_s1_begintransfer,                                          --                                                         .begintransfer
			rs232_uart_s1_chipselect                                             => mm_interconnect_2_rs232_uart_s1_chipselect,                                             --                                                         .chipselect
			rst_controller_avalon_rst_controller_slave_address                   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,                   --               rst_controller_avalon_rst_controller_slave.address
			rst_controller_avalon_rst_controller_slave_write                     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,                     --                                                         .write
			rst_controller_avalon_rst_controller_slave_read                      => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,                      --                                                         .read
			rst_controller_avalon_rst_controller_slave_readdata                  => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,                  --                                                         .readdata
			rst_controller_avalon_rst_controller_slave_writedata                 => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,                 --                                                         .writedata
			rst_controller_avalon_rst_controller_slave_waitrequest               => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest,               --                                                         .waitrequest
			rtcc_alarm_s1_address                                                => mm_interconnect_2_rtcc_alarm_s1_address,                                                --                                            rtcc_alarm_s1.address
			rtcc_alarm_s1_readdata                                               => mm_interconnect_2_rtcc_alarm_s1_readdata,                                               --                                                         .readdata
			rtcc_cs_n_s1_address                                                 => mm_interconnect_2_rtcc_cs_n_s1_address,                                                 --                                             rtcc_cs_n_s1.address
			rtcc_cs_n_s1_write                                                   => mm_interconnect_2_rtcc_cs_n_s1_write,                                                   --                                                         .write
			rtcc_cs_n_s1_readdata                                                => mm_interconnect_2_rtcc_cs_n_s1_readdata,                                                --                                                         .readdata
			rtcc_cs_n_s1_writedata                                               => mm_interconnect_2_rtcc_cs_n_s1_writedata,                                               --                                                         .writedata
			rtcc_cs_n_s1_chipselect                                              => mm_interconnect_2_rtcc_cs_n_s1_chipselect,                                              --                                                         .chipselect
			rtcc_sck_s1_address                                                  => mm_interconnect_2_rtcc_sck_s1_address,                                                  --                                              rtcc_sck_s1.address
			rtcc_sck_s1_write                                                    => mm_interconnect_2_rtcc_sck_s1_write,                                                    --                                                         .write
			rtcc_sck_s1_readdata                                                 => mm_interconnect_2_rtcc_sck_s1_readdata,                                                 --                                                         .readdata
			rtcc_sck_s1_writedata                                                => mm_interconnect_2_rtcc_sck_s1_writedata,                                                --                                                         .writedata
			rtcc_sck_s1_chipselect                                               => mm_interconnect_2_rtcc_sck_s1_chipselect,                                               --                                                         .chipselect
			rtcc_sdi_s1_address                                                  => mm_interconnect_2_rtcc_sdi_s1_address,                                                  --                                              rtcc_sdi_s1.address
			rtcc_sdi_s1_write                                                    => mm_interconnect_2_rtcc_sdi_s1_write,                                                    --                                                         .write
			rtcc_sdi_s1_readdata                                                 => mm_interconnect_2_rtcc_sdi_s1_readdata,                                                 --                                                         .readdata
			rtcc_sdi_s1_writedata                                                => mm_interconnect_2_rtcc_sdi_s1_writedata,                                                --                                                         .writedata
			rtcc_sdi_s1_chipselect                                               => mm_interconnect_2_rtcc_sdi_s1_chipselect,                                               --                                                         .chipselect
			rtcc_sdo_s1_address                                                  => mm_interconnect_2_rtcc_sdo_s1_address,                                                  --                                              rtcc_sdo_s1.address
			rtcc_sdo_s1_readdata                                                 => mm_interconnect_2_rtcc_sdo_s1_readdata,                                                 --                                                         .readdata
			sd_card_wp_n_s1_address                                              => mm_interconnect_2_sd_card_wp_n_s1_address,                                              --                                          sd_card_wp_n_s1.address
			sd_card_wp_n_s1_readdata                                             => mm_interconnect_2_sd_card_wp_n_s1_readdata,                                             --                                                         .readdata
			sync_avalon_mm_slave_address                                         => mm_interconnect_2_sync_avalon_mm_slave_address,                                         --                                     sync_avalon_mm_slave.address
			sync_avalon_mm_slave_write                                           => mm_interconnect_2_sync_avalon_mm_slave_write,                                           --                                                         .write
			sync_avalon_mm_slave_read                                            => mm_interconnect_2_sync_avalon_mm_slave_read,                                            --                                                         .read
			sync_avalon_mm_slave_readdata                                        => mm_interconnect_2_sync_avalon_mm_slave_readdata,                                        --                                                         .readdata
			sync_avalon_mm_slave_writedata                                       => mm_interconnect_2_sync_avalon_mm_slave_writedata,                                       --                                                         .writedata
			sync_avalon_mm_slave_waitrequest                                     => mm_interconnect_2_sync_avalon_mm_slave_waitrequest,                                     --                                                         .waitrequest
			temp_scl_s1_address                                                  => mm_interconnect_2_temp_scl_s1_address,                                                  --                                              temp_scl_s1.address
			temp_scl_s1_write                                                    => mm_interconnect_2_temp_scl_s1_write,                                                    --                                                         .write
			temp_scl_s1_readdata                                                 => mm_interconnect_2_temp_scl_s1_readdata,                                                 --                                                         .readdata
			temp_scl_s1_writedata                                                => mm_interconnect_2_temp_scl_s1_writedata,                                                --                                                         .writedata
			temp_scl_s1_chipselect                                               => mm_interconnect_2_temp_scl_s1_chipselect,                                               --                                                         .chipselect
			temp_sda_s1_address                                                  => mm_interconnect_2_temp_sda_s1_address,                                                  --                                              temp_sda_s1.address
			temp_sda_s1_write                                                    => mm_interconnect_2_temp_sda_s1_write,                                                    --                                                         .write
			temp_sda_s1_readdata                                                 => mm_interconnect_2_temp_sda_s1_readdata,                                                 --                                                         .readdata
			temp_sda_s1_writedata                                                => mm_interconnect_2_temp_sda_s1_writedata,                                                --                                                         .writedata
			temp_sda_s1_chipselect                                               => mm_interconnect_2_temp_sda_s1_chipselect,                                               --                                                         .chipselect
			timer_1ms_s1_address                                                 => mm_interconnect_2_timer_1ms_s1_address,                                                 --                                             timer_1ms_s1.address
			timer_1ms_s1_write                                                   => mm_interconnect_2_timer_1ms_s1_write,                                                   --                                                         .write
			timer_1ms_s1_readdata                                                => mm_interconnect_2_timer_1ms_s1_readdata,                                                --                                                         .readdata
			timer_1ms_s1_writedata                                               => mm_interconnect_2_timer_1ms_s1_writedata,                                               --                                                         .writedata
			timer_1ms_s1_chipselect                                              => mm_interconnect_2_timer_1ms_s1_chipselect,                                              --                                                         .chipselect
			timer_1us_s1_address                                                 => mm_interconnect_2_timer_1us_s1_address,                                                 --                                             timer_1us_s1.address
			timer_1us_s1_write                                                   => mm_interconnect_2_timer_1us_s1_write,                                                   --                                                         .write
			timer_1us_s1_readdata                                                => mm_interconnect_2_timer_1us_s1_readdata,                                                --                                                         .readdata
			timer_1us_s1_writedata                                               => mm_interconnect_2_timer_1us_s1_writedata,                                               --                                                         .writedata
			timer_1us_s1_chipselect                                              => mm_interconnect_2_timer_1us_s1_chipselect                                               --                                                         .chipselect
		);

	mm_interconnect_3 : component MebX_Qsys_Project_mm_interconnect_3
		port map (
			m1_ddr2_memory_afi_clk_clk                                      => m1_ddr2_memory_afi_clk_clk,                              --                                    m1_ddr2_memory_afi_clk.clk
			m1_ddr2_memory_afi_half_clk_clk                                 => m1_ddr2_memory_afi_half_clk_clk,                         --                               m1_ddr2_memory_afi_half_clk.clk
			m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset            => rst_controller_005_reset_out_reset,                      --            m1_clock_bridge_m0_reset_reset_bridge_in_reset.reset
			m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset => rst_controller_008_reset_out_reset,                      -- m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
			m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           => rst_controller_008_reset_out_reset,                      --           m1_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
			m1_clock_bridge_m0_address                                      => m1_clock_bridge_m0_address,                              --                                        m1_clock_bridge_m0.address
			m1_clock_bridge_m0_waitrequest                                  => m1_clock_bridge_m0_waitrequest,                          --                                                          .waitrequest
			m1_clock_bridge_m0_burstcount                                   => m1_clock_bridge_m0_burstcount,                           --                                                          .burstcount
			m1_clock_bridge_m0_byteenable                                   => m1_clock_bridge_m0_byteenable,                           --                                                          .byteenable
			m1_clock_bridge_m0_read                                         => m1_clock_bridge_m0_read,                                 --                                                          .read
			m1_clock_bridge_m0_readdata                                     => m1_clock_bridge_m0_readdata,                             --                                                          .readdata
			m1_clock_bridge_m0_readdatavalid                                => m1_clock_bridge_m0_readdatavalid,                        --                                                          .readdatavalid
			m1_clock_bridge_m0_write                                        => m1_clock_bridge_m0_write,                                --                                                          .write
			m1_clock_bridge_m0_writedata                                    => m1_clock_bridge_m0_writedata,                            --                                                          .writedata
			m1_clock_bridge_m0_debugaccess                                  => m1_clock_bridge_m0_debugaccess,                          --                                                          .debugaccess
			m1_ddr2_memory_avl_address                                      => mm_interconnect_3_m1_ddr2_memory_avl_address,            --                                        m1_ddr2_memory_avl.address
			m1_ddr2_memory_avl_write                                        => mm_interconnect_3_m1_ddr2_memory_avl_write,              --                                                          .write
			m1_ddr2_memory_avl_read                                         => mm_interconnect_3_m1_ddr2_memory_avl_read,               --                                                          .read
			m1_ddr2_memory_avl_readdata                                     => mm_interconnect_3_m1_ddr2_memory_avl_readdata,           --                                                          .readdata
			m1_ddr2_memory_avl_writedata                                    => mm_interconnect_3_m1_ddr2_memory_avl_writedata,          --                                                          .writedata
			m1_ddr2_memory_avl_beginbursttransfer                           => mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer, --                                                          .beginbursttransfer
			m1_ddr2_memory_avl_burstcount                                   => mm_interconnect_3_m1_ddr2_memory_avl_burstcount,         --                                                          .burstcount
			m1_ddr2_memory_avl_byteenable                                   => mm_interconnect_3_m1_ddr2_memory_avl_byteenable,         --                                                          .byteenable
			m1_ddr2_memory_avl_readdatavalid                                => mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid,      --                                                          .readdatavalid
			m1_ddr2_memory_avl_waitrequest                                  => mm_interconnect_3_m1_ddr2_memory_avl_inv                 --                                                          .waitrequest
		);

	irq_mapper : component MebX_Qsys_Project_irq_mapper
		port map (
			clk            => m2_ddr2_memory_afi_half_clk_clk,    --        clk.clk
			reset          => rst_controller_006_reset_out_reset, --  clk_reset.reset
			receiver0_irq  => irq_mapper_receiver0_irq,           --  receiver0.irq
			receiver1_irq  => irq_mapper_receiver1_irq,           --  receiver1.irq
			receiver2_irq  => irq_mapper_receiver2_irq,           --  receiver2.irq
			receiver3_irq  => irq_mapper_receiver3_irq,           --  receiver3.irq
			receiver4_irq  => irq_mapper_receiver4_irq,           --  receiver4.irq
			receiver5_irq  => irq_mapper_receiver5_irq,           --  receiver5.irq
			receiver6_irq  => irq_mapper_receiver6_irq,           --  receiver6.irq
			receiver7_irq  => irq_mapper_receiver7_irq,           --  receiver7.irq
			receiver8_irq  => irq_mapper_receiver8_irq,           --  receiver8.irq
			receiver9_irq  => irq_mapper_receiver9_irq,           --  receiver9.irq
			receiver10_irq => irq_mapper_receiver10_irq,          -- receiver10.irq
			receiver11_irq => irq_mapper_receiver11_irq,          -- receiver11.irq
			receiver12_irq => irq_mapper_receiver12_irq,          -- receiver12.irq
			receiver13_irq => irq_mapper_receiver13_irq,          -- receiver13.irq
			receiver14_irq => irq_mapper_receiver14_irq,          -- receiver14.irq
			receiver15_irq => irq_mapper_receiver15_irq,          -- receiver15.irq
			sender_irq     => nios2_gen2_0_irq_irq                --     sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_006_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver5_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_006_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver6_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_007_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_006_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver7_irq            --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_006_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver8_irq            --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_006_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver14_irq           --             sender.irq
		);

	rst_controller_001 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => clk50_clk,                          --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component mebx_qsys_project_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component mebx_qsys_project_rst_controller_004
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => rst_reset_n_ports_inv,              -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,    --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_005 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m1_ddr2_memory_afi_half_clk_clk,    --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_006 : component mebx_qsys_project_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_006_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_007 : component mebx_qsys_project_rst_controller_004
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                   -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_rs232_reset, -- reset_in1.reset
			clk            => clk50_clk,                               --       clk.clk
			reset_out      => rst_controller_007_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                    -- (terminated)
			reset_req_in0  => '0',                                     -- (terminated)
			reset_req_in1  => '0',                                     -- (terminated)
			reset_in2      => '0',                                     -- (terminated)
			reset_req_in2  => '0',                                     -- (terminated)
			reset_in3      => '0',                                     -- (terminated)
			reset_req_in3  => '0',                                     -- (terminated)
			reset_in4      => '0',                                     -- (terminated)
			reset_req_in4  => '0',                                     -- (terminated)
			reset_in5      => '0',                                     -- (terminated)
			reset_req_in5  => '0',                                     -- (terminated)
			reset_in6      => '0',                                     -- (terminated)
			reset_req_in6  => '0',                                     -- (terminated)
			reset_in7      => '0',                                     -- (terminated)
			reset_req_in7  => '0',                                     -- (terminated)
			reset_in8      => '0',                                     -- (terminated)
			reset_req_in8  => '0',                                     -- (terminated)
			reset_in9      => '0',                                     -- (terminated)
			reset_req_in9  => '0',                                     -- (terminated)
			reset_in10     => '0',                                     -- (terminated)
			reset_req_in10 => '0',                                     -- (terminated)
			reset_in11     => '0',                                     -- (terminated)
			reset_req_in11 => '0',                                     -- (terminated)
			reset_in12     => '0',                                     -- (terminated)
			reset_req_in12 => '0',                                     -- (terminated)
			reset_in13     => '0',                                     -- (terminated)
			reset_req_in13 => '0',                                     -- (terminated)
			reset_in14     => '0',                                     -- (terminated)
			reset_req_in14 => '0',                                     -- (terminated)
			reset_in15     => '0',                                     -- (terminated)
			reset_req_in15 => '0'                                      -- (terminated)
		);

	rst_controller_008 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m1_ddr2_memory_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_008_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_reset_n_ports_inv <= not rst_reset_n;

	mm_interconnect_0_m2_ddr2_memory_avl_inv <= not m2_ddr2_memory_avl_waitrequest;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv <= not mm_interconnect_2_m1_ddr2_i2c_sda_s1_write;

	mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv <= not mm_interconnect_2_m1_ddr2_i2c_scl_s1_write;

	mm_interconnect_2_pio_led_s1_write_ports_inv <= not mm_interconnect_2_pio_led_s1_write;

	mm_interconnect_2_timer_1ms_s1_write_ports_inv <= not mm_interconnect_2_timer_1ms_s1_write;

	mm_interconnect_2_timer_1us_s1_write_ports_inv <= not mm_interconnect_2_timer_1us_s1_write;

	mm_interconnect_2_temp_scl_s1_write_ports_inv <= not mm_interconnect_2_temp_scl_s1_write;

	mm_interconnect_2_temp_sda_s1_write_ports_inv <= not mm_interconnect_2_temp_sda_s1_write;

	mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv <= not mm_interconnect_2_m2_ddr2_i2c_sda_s1_write;

	mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv <= not mm_interconnect_2_m2_ddr2_i2c_scl_s1_write;

	mm_interconnect_2_csense_sdi_s1_write_ports_inv <= not mm_interconnect_2_csense_sdi_s1_write;

	mm_interconnect_2_csense_sck_s1_write_ports_inv <= not mm_interconnect_2_csense_sck_s1_write;

	mm_interconnect_2_csense_cs_n_s1_write_ports_inv <= not mm_interconnect_2_csense_cs_n_s1_write;

	mm_interconnect_2_csense_adc_fo_s1_write_ports_inv <= not mm_interconnect_2_csense_adc_fo_s1_write;

	mm_interconnect_2_pio_led_painel_s1_write_ports_inv <= not mm_interconnect_2_pio_led_painel_s1_write;

	mm_interconnect_2_rtcc_sdi_s1_write_ports_inv <= not mm_interconnect_2_rtcc_sdi_s1_write;

	mm_interconnect_2_rtcc_sck_s1_write_ports_inv <= not mm_interconnect_2_rtcc_sck_s1_write;

	mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv <= not mm_interconnect_2_rtcc_cs_n_s1_write;

	mm_interconnect_2_rs232_uart_s1_read_ports_inv <= not mm_interconnect_2_rs232_uart_s1_read;

	mm_interconnect_2_rs232_uart_s1_write_ports_inv <= not mm_interconnect_2_rs232_uart_s1_write;

	mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv <= not mm_interconnect_2_pio_ctrl_io_lvds_s1_write;

	mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write_ports_inv <= not mm_interconnect_2_pio_spw_demux_ch_1_select_s1_write;

	mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write_ports_inv <= not mm_interconnect_2_pio_spw_demux_ch_2_select_s1_write;

	mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write_ports_inv <= not mm_interconnect_2_pio_spw_demux_ch_3_select_s1_write;

	mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write_ports_inv <= not mm_interconnect_2_pio_spw_demux_ch_4_select_s1_write;

	mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write_ports_inv <= not mm_interconnect_2_pio_ftdi_umft601a_module_reset_s1_write;

	mm_interconnect_2_pio_iso_logic_signal_enable_s1_write_ports_inv <= not mm_interconnect_2_pio_iso_logic_signal_enable_s1_write;

	mm_interconnect_3_m1_ddr2_memory_avl_inv <= not m1_ddr2_memory_avl_waitrequest;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_006_reset_out_reset_ports_inv <= not rst_controller_006_reset_out_reset;

	rst_controller_007_reset_out_reset_ports_inv <= not rst_controller_007_reset_out_reset;

end architecture rtl; -- of MebX_Qsys_Project
